-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Oct 8 2022 16:56:32

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "LED_blink" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of LED_blink
entity LED_blink is
port (
    o_LED_3 : out std_logic;
    o_LED_1 : out std_logic;
    i_Clk : in std_logic;
    o_LED_4 : out std_logic;
    o_LED_2 : out std_logic);
end LED_blink;

-- Architecture of LED_blink
-- View name is \INTERFACE\
architecture \INTERFACE\ of LED_blink is

signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \o_LED_33_0\ : std_logic;
signal \o_LED_33_1\ : std_logic;
signal \o_LED_33_2\ : std_logic;
signal \o_LED_33_3\ : std_logic;
signal \o_LED_33_4\ : std_logic;
signal \o_LED_33_5\ : std_logic;
signal \o_LED_33_6\ : std_logic;
signal \o_LED_33\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \o_LED_33_THRU_CO_cascade_\ : std_logic;
signal \o_LED_3_c\ : std_logic;
signal \o_LED_33_2_and\ : std_logic;
signal \o_LED_33_1_and\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \o_LED_23_0\ : std_logic;
signal \o_LED_23_1\ : std_logic;
signal \o_LED_23_2\ : std_logic;
signal \o_LED_23_3\ : std_logic;
signal \o_LED_23_4\ : std_logic;
signal \o_LED_23_5\ : std_logic;
signal \o_LED_23_6\ : std_logic;
signal \o_LED_23\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \o_LED_33_4_and\ : std_logic;
signal \o_LED_33_3_and\ : std_logic;
signal \o_LED_33_5_and\ : std_logic;
signal \o_LED_33_0_and\ : std_logic;
signal \o_LED_33_6_and\ : std_logic;
signal \o_LED_33_THRU_CO\ : std_logic;
signal \o_LED_33_7_and\ : std_logic;
signal \o_LED_23_2_and\ : std_logic;
signal \o_LED_23_3_and\ : std_logic;
signal \o_LED_23_1_and\ : std_logic;
signal \o_LED_23_0_and\ : std_logic;
signal \o_LED_23_7_and\ : std_logic;
signal \o_LED_23_5_and\ : std_logic;
signal \o_LED_2_c\ : std_logic;
signal \o_LED_23_6_and\ : std_logic;
signal \o_LED_23_4_and\ : std_logic;
signal \o_LED_23_THRU_CO\ : std_logic;
signal \r_count_2hzZ0Z_0\ : std_logic;
signal \r_count_2hzZ0Z_1\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \r_count_2hzZ0Z_2\ : std_logic;
signal un2_r_count_2hz_1_cry_1 : std_logic;
signal \r_count_2hzZ0Z_3\ : std_logic;
signal un2_r_count_2hz_1_cry_2 : std_logic;
signal \r_count_2hzZ0Z_4\ : std_logic;
signal \un2_r_count_2hz_1_cry_3_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_3 : std_logic;
signal \r_count_2hzZ0Z_5\ : std_logic;
signal un2_r_count_2hz_1_cry_4 : std_logic;
signal \r_count_2hzZ0Z_6\ : std_logic;
signal un2_r_count_2hz_1_cry_5 : std_logic;
signal \r_count_2hzZ0Z_7\ : std_logic;
signal un2_r_count_2hz_1_cry_6 : std_logic;
signal \r_count_2hzZ0Z_8\ : std_logic;
signal un2_r_count_2hz_1_cry_7 : std_logic;
signal un2_r_count_2hz_1_cry_8 : std_logic;
signal \r_count_2hzZ0Z_9\ : std_logic;
signal \un2_r_count_2hz_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \r_count_2hzZ0Z_10\ : std_logic;
signal \un2_r_count_2hz_1_cry_9_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_9 : std_logic;
signal \r_count_2hzZ0Z_11\ : std_logic;
signal \un2_r_count_2hz_1_cry_10_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_10 : std_logic;
signal \r_count_2hzZ0Z_12\ : std_logic;
signal \un2_r_count_2hz_1_cry_11_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_11 : std_logic;
signal \r_count_2hzZ0Z_13\ : std_logic;
signal un2_r_count_2hz_1_cry_12 : std_logic;
signal \r_count_2hzZ0Z_14\ : std_logic;
signal \un2_r_count_2hz_1_cry_13_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_13 : std_logic;
signal \r_count_2hzZ0Z_15\ : std_logic;
signal un2_r_count_2hz_1_cry_14 : std_logic;
signal \r_count_2hzZ0Z_16\ : std_logic;
signal \un2_r_count_2hz_1_cry_15_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_15 : std_logic;
signal un2_r_count_2hz_1_cry_16 : std_logic;
signal \r_count_2hzZ0Z_17\ : std_logic;
signal \un2_r_count_2hz_1_cry_16_THRU_CO\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \r_count_2hzZ0Z_18\ : std_logic;
signal \un2_r_count_2hz_1_cry_17_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_17 : std_logic;
signal \r_count_2hzZ0Z_19\ : std_logic;
signal \un2_r_count_2hz_1_cry_18_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_18 : std_logic;
signal \r_count_2hzZ0Z_20\ : std_logic;
signal \un2_r_count_2hz_1_cry_19_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_19 : std_logic;
signal \r_count_2hzZ0Z_21\ : std_logic;
signal un2_r_count_2hz_1_cry_20 : std_logic;
signal \r_count_2hzZ0Z_22\ : std_logic;
signal \un2_r_count_2hz_1_cry_21_THRU_CO\ : std_logic;
signal un2_r_count_2hz_1_cry_21 : std_logic;
signal \r_count_2hzZ0Z_23\ : std_logic;
signal un2_r_count_2hz_1_cry_22 : std_logic;
signal \r_count_2hzZ0Z_24\ : std_logic;
signal un2_r_count_2hz_1_cry_23 : std_logic;
signal un2_r_count_2hz_1_cry_24 : std_logic;
signal \r_count_2hzZ0Z_25\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \r_count_2hzZ0Z_26\ : std_logic;
signal un2_r_count_2hz_1_cry_25 : std_logic;
signal \r_count_2hzZ0Z_27\ : std_logic;
signal un2_r_count_2hz_1_cry_26 : std_logic;
signal \r_count_2hzZ0Z_28\ : std_logic;
signal un2_r_count_2hz_1_cry_27 : std_logic;
signal \r_count_2hzZ0Z_29\ : std_logic;
signal un2_r_count_2hz_1_cry_28 : std_logic;
signal \r_count_2hzZ0Z_30\ : std_logic;
signal un2_r_count_2hz_1_cry_29 : std_logic;
signal un2_r_count_2hz_1_cry_30 : std_logic;
signal \r_count_2hzZ0Z_31\ : std_logic;
signal \o_LED_4_c\ : std_logic;
signal \r_count_5hzZ0Z_0\ : std_logic;
signal \r_count_5hzZ0Z_1\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \r_count_5hzZ0Z_2\ : std_logic;
signal un2_r_count_5hz_1_cry_1 : std_logic;
signal \r_count_5hzZ0Z_3\ : std_logic;
signal un2_r_count_5hz_1_cry_2 : std_logic;
signal \r_count_5hzZ0Z_4\ : std_logic;
signal \un2_r_count_5hz_1_cry_3_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_3 : std_logic;
signal \r_count_5hzZ0Z_5\ : std_logic;
signal un2_r_count_5hz_1_cry_4 : std_logic;
signal \r_count_5hzZ0Z_6\ : std_logic;
signal un2_r_count_5hz_1_cry_5 : std_logic;
signal \r_count_5hzZ0Z_7\ : std_logic;
signal \un2_r_count_5hz_1_cry_6_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_6 : std_logic;
signal \r_count_5hzZ0Z_8\ : std_logic;
signal un2_r_count_5hz_1_cry_7 : std_logic;
signal un2_r_count_5hz_1_cry_8 : std_logic;
signal \r_count_5hzZ0Z_9\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \r_count_5hzZ0Z_10\ : std_logic;
signal un2_r_count_5hz_1_cry_9 : std_logic;
signal \r_count_5hzZ0Z_11\ : std_logic;
signal un2_r_count_5hz_1_cry_10 : std_logic;
signal \r_count_5hzZ0Z_12\ : std_logic;
signal \un2_r_count_5hz_1_cry_11_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_11 : std_logic;
signal \r_count_5hzZ0Z_13\ : std_logic;
signal un2_r_count_5hz_1_cry_12 : std_logic;
signal \r_count_5hzZ0Z_14\ : std_logic;
signal \un2_r_count_5hz_1_cry_13_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_13 : std_logic;
signal \r_count_5hzZ0Z_15\ : std_logic;
signal \un2_r_count_5hz_1_cry_14_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_14 : std_logic;
signal \r_count_5hzZ0Z_16\ : std_logic;
signal \un2_r_count_5hz_1_cry_15_THRU_CO\ : std_logic;
signal un2_r_count_5hz_1_cry_15 : std_logic;
signal un2_r_count_5hz_1_cry_16 : std_logic;
signal \r_count_5hzZ0Z_17\ : std_logic;
signal \un2_r_count_5hz_1_cry_16_THRU_CO\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \r_count_5hzZ0Z_18\ : std_logic;
signal un2_r_count_5hz_1_cry_17 : std_logic;
signal \r_count_5hzZ0Z_19\ : std_logic;
signal un2_r_count_5hz_1_cry_18 : std_logic;
signal \r_count_5hzZ0Z_20\ : std_logic;
signal un2_r_count_5hz_1_cry_19 : std_logic;
signal \r_count_5hzZ0Z_21\ : std_logic;
signal un2_r_count_5hz_1_cry_20 : std_logic;
signal \r_count_5hzZ0Z_22\ : std_logic;
signal un2_r_count_5hz_1_cry_21 : std_logic;
signal \r_count_5hzZ0Z_23\ : std_logic;
signal un2_r_count_5hz_1_cry_22 : std_logic;
signal \r_count_5hzZ0Z_24\ : std_logic;
signal un2_r_count_5hz_1_cry_23 : std_logic;
signal un2_r_count_5hz_1_cry_24 : std_logic;
signal \r_count_5hzZ0Z_25\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \r_count_5hzZ0Z_26\ : std_logic;
signal un2_r_count_5hz_1_cry_25 : std_logic;
signal \r_count_5hzZ0Z_27\ : std_logic;
signal un2_r_count_5hz_1_cry_26 : std_logic;
signal \r_count_5hzZ0Z_28\ : std_logic;
signal un2_r_count_5hz_1_cry_27 : std_logic;
signal \r_count_5hzZ0Z_29\ : std_logic;
signal un2_r_count_5hz_1_cry_28 : std_logic;
signal \r_count_5hzZ0Z_30\ : std_logic;
signal un2_r_count_5hz_1_cry_29 : std_logic;
signal un2_r_count_5hz_1_cry_30 : std_logic;
signal \r_count_5hzZ0Z_31\ : std_logic;
signal \o_LED_43_0_and\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \o_LED_43_0\ : std_logic;
signal \o_LED_43_1\ : std_logic;
signal \o_LED_43_3_and\ : std_logic;
signal \o_LED_43_2\ : std_logic;
signal \o_LED_43_3\ : std_logic;
signal \o_LED_43_4\ : std_logic;
signal \o_LED_43_5\ : std_logic;
signal \o_LED_43_6\ : std_logic;
signal \o_LED_43\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \o_LED_43_THRU_CO_cascade_\ : std_logic;
signal \o_LED_43_1_and\ : std_logic;
signal \o_LED_43_2_and\ : std_logic;
signal \o_LED_43_THRU_CO\ : std_logic;
signal \bfn_11_1_0_\ : std_logic;
signal \o_LED_13_0\ : std_logic;
signal \o_LED_13_1\ : std_logic;
signal \o_LED_13_2\ : std_logic;
signal \o_LED_13_3\ : std_logic;
signal \o_LED_13_4\ : std_logic;
signal \o_LED_13_5\ : std_logic;
signal \o_LED_13_6\ : std_logic;
signal \o_LED_13\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \o_LED_13_THRU_CO_cascade_\ : std_logic;
signal \o_LED_13_1_and\ : std_logic;
signal \o_LED_1_c\ : std_logic;
signal \o_LED_13_4_and\ : std_logic;
signal \o_LED_13_5_and\ : std_logic;
signal \o_LED_13_6_and\ : std_logic;
signal \o_LED_13_7_and\ : std_logic;
signal \o_LED_43_4_and\ : std_logic;
signal \r_count_1hzZ0Z_0\ : std_logic;
signal \r_count_1hzZ0Z_1\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \r_count_1hzZ0Z_2\ : std_logic;
signal un2_r_count_1hz_1_cry_1 : std_logic;
signal \r_count_1hzZ0Z_3\ : std_logic;
signal un2_r_count_1hz_1_cry_2 : std_logic;
signal \r_count_1hzZ0Z_4\ : std_logic;
signal un2_r_count_1hz_1_cry_3 : std_logic;
signal \r_count_1hzZ0Z_5\ : std_logic;
signal \un2_r_count_1hz_1_cry_4_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_4 : std_logic;
signal \r_count_1hzZ0Z_6\ : std_logic;
signal un2_r_count_1hz_1_cry_5 : std_logic;
signal \r_count_1hzZ0Z_7\ : std_logic;
signal un2_r_count_1hz_1_cry_6 : std_logic;
signal \r_count_1hzZ0Z_8\ : std_logic;
signal un2_r_count_1hz_1_cry_7 : std_logic;
signal un2_r_count_1hz_1_cry_8 : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \r_count_1hzZ0Z_10\ : std_logic;
signal \un2_r_count_1hz_1_cry_9_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_9 : std_logic;
signal \r_count_1hzZ0Z_11\ : std_logic;
signal \un2_r_count_1hz_1_cry_10_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_10 : std_logic;
signal \r_count_1hzZ0Z_12\ : std_logic;
signal \un2_r_count_1hz_1_cry_11_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_11 : std_logic;
signal \r_count_1hzZ0Z_13\ : std_logic;
signal \un2_r_count_1hz_1_cry_12_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_12 : std_logic;
signal un2_r_count_1hz_1_cry_13 : std_logic;
signal \r_count_1hzZ0Z_15\ : std_logic;
signal \un2_r_count_1hz_1_cry_14_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_14 : std_logic;
signal un2_r_count_1hz_1_cry_15 : std_logic;
signal un2_r_count_1hz_1_cry_16 : std_logic;
signal \r_count_1hzZ0Z_17\ : std_logic;
signal \un2_r_count_1hz_1_cry_16_THRU_CO\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \r_count_1hzZ0Z_18\ : std_logic;
signal \un2_r_count_1hz_1_cry_17_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_17 : std_logic;
signal \r_count_1hzZ0Z_19\ : std_logic;
signal \un2_r_count_1hz_1_cry_18_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_18 : std_logic;
signal \r_count_1hzZ0Z_20\ : std_logic;
signal \un2_r_count_1hz_1_cry_19_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_19 : std_logic;
signal \r_count_1hzZ0Z_21\ : std_logic;
signal \un2_r_count_1hz_1_cry_20_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_20 : std_logic;
signal un2_r_count_1hz_1_cry_21 : std_logic;
signal \r_count_1hzZ0Z_23\ : std_logic;
signal \un2_r_count_1hz_1_cry_22_THRU_CO\ : std_logic;
signal un2_r_count_1hz_1_cry_22 : std_logic;
signal un2_r_count_1hz_1_cry_23 : std_logic;
signal un2_r_count_1hz_1_cry_24 : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal un2_r_count_1hz_1_cry_25 : std_logic;
signal un2_r_count_1hz_1_cry_26 : std_logic;
signal un2_r_count_1hz_1_cry_27 : std_logic;
signal un2_r_count_1hz_1_cry_28 : std_logic;
signal un2_r_count_1hz_1_cry_29 : std_logic;
signal un2_r_count_1hz_1_cry_30 : std_logic;
signal \r_count_1hzZ0Z_29\ : std_logic;
signal \r_count_1hzZ0Z_31\ : std_logic;
signal \r_count_1hzZ0Z_28\ : std_logic;
signal \r_count_1hzZ0Z_30\ : std_logic;
signal \o_LED_43_7_and\ : std_logic;
signal \o_LED_13_THRU_CO\ : std_logic;
signal \o_LED_13_0_and\ : std_logic;
signal \o_LED_13_3_and\ : std_logic;
signal \o_LED_13_2_and\ : std_logic;
signal \r_count_10hzZ0Z_0\ : std_logic;
signal \r_count_10hzZ0Z_1\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \r_count_10hzZ0Z_2\ : std_logic;
signal un2_r_count_10hz_1_cry_1 : std_logic;
signal \r_count_10hzZ0Z_3\ : std_logic;
signal un2_r_count_10hz_1_cry_2 : std_logic;
signal \r_count_10hzZ0Z_4\ : std_logic;
signal \un2_r_count_10hz_1_cry_3_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_3 : std_logic;
signal \r_count_10hzZ0Z_5\ : std_logic;
signal un2_r_count_10hz_1_cry_4 : std_logic;
signal \r_count_10hzZ0Z_6\ : std_logic;
signal \un2_r_count_10hz_1_cry_5_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_5 : std_logic;
signal \r_count_10hzZ0Z_7\ : std_logic;
signal \un2_r_count_10hz_1_cry_6_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_6 : std_logic;
signal \r_count_10hzZ0Z_8\ : std_logic;
signal un2_r_count_10hz_1_cry_7 : std_logic;
signal un2_r_count_10hz_1_cry_8 : std_logic;
signal \r_count_10hzZ0Z_9\ : std_logic;
signal \un2_r_count_10hz_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \r_count_10hzZ0Z_10\ : std_logic;
signal un2_r_count_10hz_1_cry_9 : std_logic;
signal \r_count_10hzZ0Z_11\ : std_logic;
signal un2_r_count_10hz_1_cry_10 : std_logic;
signal \r_count_10hzZ0Z_12\ : std_logic;
signal \un2_r_count_10hz_1_cry_11_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_11 : std_logic;
signal \r_count_10hzZ0Z_13\ : std_logic;
signal un2_r_count_10hz_1_cry_12 : std_logic;
signal \r_count_10hzZ0Z_14\ : std_logic;
signal un2_r_count_10hz_1_cry_13 : std_logic;
signal \r_count_10hzZ0Z_15\ : std_logic;
signal un2_r_count_10hz_1_cry_14 : std_logic;
signal \r_count_10hzZ0Z_16\ : std_logic;
signal \un2_r_count_10hz_1_cry_15_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_15 : std_logic;
signal un2_r_count_10hz_1_cry_16 : std_logic;
signal \r_count_10hzZ0Z_17\ : std_logic;
signal \un2_r_count_10hz_1_cry_16_THRU_CO\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \r_count_10hzZ0Z_18\ : std_logic;
signal un2_r_count_10hz_1_cry_17 : std_logic;
signal \r_count_10hzZ0Z_19\ : std_logic;
signal un2_r_count_10hz_1_cry_18 : std_logic;
signal \r_count_10hzZ0Z_20\ : std_logic;
signal \un2_r_count_10hz_1_cry_19_THRU_CO\ : std_logic;
signal un2_r_count_10hz_1_cry_19 : std_logic;
signal \r_count_10hzZ0Z_21\ : std_logic;
signal un2_r_count_10hz_1_cry_20 : std_logic;
signal \r_count_10hzZ0Z_22\ : std_logic;
signal un2_r_count_10hz_1_cry_21 : std_logic;
signal \r_count_10hzZ0Z_23\ : std_logic;
signal un2_r_count_10hz_1_cry_22 : std_logic;
signal \r_count_10hzZ0Z_24\ : std_logic;
signal un2_r_count_10hz_1_cry_23 : std_logic;
signal un2_r_count_10hz_1_cry_24 : std_logic;
signal \r_count_10hzZ0Z_25\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \r_count_10hzZ0Z_26\ : std_logic;
signal un2_r_count_10hz_1_cry_25 : std_logic;
signal \r_count_10hzZ0Z_27\ : std_logic;
signal un2_r_count_10hz_1_cry_26 : std_logic;
signal \r_count_10hzZ0Z_28\ : std_logic;
signal un2_r_count_10hz_1_cry_27 : std_logic;
signal \r_count_10hzZ0Z_29\ : std_logic;
signal un2_r_count_10hz_1_cry_28 : std_logic;
signal \r_count_10hzZ0Z_30\ : std_logic;
signal un2_r_count_10hz_1_cry_29 : std_logic;
signal un2_r_count_10hz_1_cry_30 : std_logic;
signal \r_count_10hzZ0Z_31\ : std_logic;
signal \i_Clk_c_g\ : std_logic;
signal \r_count_1hzZ0Z_14\ : std_logic;
signal \r_count_1hzZ0Z_22\ : std_logic;
signal \r_count_1hzZ0Z_9\ : std_logic;
signal \r_count_1hzZ0Z_16\ : std_logic;
signal \o_LED_43_5_and\ : std_logic;
signal \r_count_1hzZ0Z_25\ : std_logic;
signal \r_count_1hzZ0Z_26\ : std_logic;
signal \r_count_1hzZ0Z_24\ : std_logic;
signal \r_count_1hzZ0Z_27\ : std_logic;
signal \o_LED_43_6_and\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \i_Clk_wire\ : std_logic;
signal \o_LED_1_wire\ : std_logic;
signal \o_LED_2_wire\ : std_logic;
signal \o_LED_4_wire\ : std_logic;
signal \o_LED_3_wire\ : std_logic;

begin
    \i_Clk_wire\ <= i_Clk;
    o_LED_1 <= \o_LED_1_wire\;
    o_LED_2 <= \o_LED_2_wire\;
    o_LED_4 <= \o_LED_4_wire\;
    o_LED_3 <= \o_LED_3_wire\;

    \i_Clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6647\,
            GLOBALBUFFEROUTPUT => \i_Clk_c_g\
        );

    \i_Clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6649\,
            DIN => \N__6648\,
            DOUT => \N__6647\,
            PACKAGEPIN => \i_Clk_wire\
        );

    \i_Clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6649\,
            PADOUT => \N__6648\,
            PADIN => \N__6647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6638\,
            DIN => \N__6637\,
            DOUT => \N__6636\,
            PACKAGEPIN => \o_LED_1_wire\
        );

    \o_LED_1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6638\,
            PADOUT => \N__6637\,
            PADIN => \N__6636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6629\,
            DIN => \N__6628\,
            DOUT => \N__6627\,
            PACKAGEPIN => \o_LED_2_wire\
        );

    \o_LED_2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6629\,
            PADOUT => \N__6628\,
            PADIN => \N__6627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3376\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6620\,
            DIN => \N__6619\,
            DOUT => \N__6618\,
            PACKAGEPIN => \o_LED_4_wire\
        );

    \o_LED_4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6620\,
            PADOUT => \N__6619\,
            PADIN => \N__6618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_LED_3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6611\,
            DIN => \N__6610\,
            DOUT => \N__6609\,
            PACKAGEPIN => \o_LED_3_wire\
        );

    \o_LED_3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6611\,
            PADOUT => \N__6610\,
            PADIN => \N__6609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3208\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1415\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6588\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6585\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6588\,
            I => \r_count_10hzZ0Z_27\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6585\,
            I => \r_count_10hzZ0Z_27\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6580\,
            I => un2_r_count_10hz_1_cry_26
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__6577\,
            I => \N__6573\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6570\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6567\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6570\,
            I => \r_count_10hzZ0Z_28\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6567\,
            I => \r_count_10hzZ0Z_28\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6562\,
            I => un2_r_count_10hz_1_cry_27
        );

    \I__1404\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6555\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6552\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6555\,
            I => \r_count_10hzZ0Z_29\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6552\,
            I => \r_count_10hzZ0Z_29\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6547\,
            I => un2_r_count_10hz_1_cry_28
        );

    \I__1399\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6540\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6537\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6540\,
            I => \r_count_10hzZ0Z_30\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6537\,
            I => \r_count_10hzZ0Z_30\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6532\,
            I => un2_r_count_10hz_1_cry_29
        );

    \I__1394\ : InMux
    port map (
            O => \N__6529\,
            I => un2_r_count_10hz_1_cry_30
        );

    \I__1393\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6522\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6519\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6522\,
            I => \r_count_10hzZ0Z_31\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6519\,
            I => \r_count_10hzZ0Z_31\
        );

    \I__1389\ : ClkMux
    port map (
            O => \N__6514\,
            I => \N__6421\
        );

    \I__1388\ : ClkMux
    port map (
            O => \N__6513\,
            I => \N__6421\
        );

    \I__1387\ : ClkMux
    port map (
            O => \N__6512\,
            I => \N__6421\
        );

    \I__1386\ : ClkMux
    port map (
            O => \N__6511\,
            I => \N__6421\
        );

    \I__1385\ : ClkMux
    port map (
            O => \N__6510\,
            I => \N__6421\
        );

    \I__1384\ : ClkMux
    port map (
            O => \N__6509\,
            I => \N__6421\
        );

    \I__1383\ : ClkMux
    port map (
            O => \N__6508\,
            I => \N__6421\
        );

    \I__1382\ : ClkMux
    port map (
            O => \N__6507\,
            I => \N__6421\
        );

    \I__1381\ : ClkMux
    port map (
            O => \N__6506\,
            I => \N__6421\
        );

    \I__1380\ : ClkMux
    port map (
            O => \N__6505\,
            I => \N__6421\
        );

    \I__1379\ : ClkMux
    port map (
            O => \N__6504\,
            I => \N__6421\
        );

    \I__1378\ : ClkMux
    port map (
            O => \N__6503\,
            I => \N__6421\
        );

    \I__1377\ : ClkMux
    port map (
            O => \N__6502\,
            I => \N__6421\
        );

    \I__1376\ : ClkMux
    port map (
            O => \N__6501\,
            I => \N__6421\
        );

    \I__1375\ : ClkMux
    port map (
            O => \N__6500\,
            I => \N__6421\
        );

    \I__1374\ : ClkMux
    port map (
            O => \N__6499\,
            I => \N__6421\
        );

    \I__1373\ : ClkMux
    port map (
            O => \N__6498\,
            I => \N__6421\
        );

    \I__1372\ : ClkMux
    port map (
            O => \N__6497\,
            I => \N__6421\
        );

    \I__1371\ : ClkMux
    port map (
            O => \N__6496\,
            I => \N__6421\
        );

    \I__1370\ : ClkMux
    port map (
            O => \N__6495\,
            I => \N__6421\
        );

    \I__1369\ : ClkMux
    port map (
            O => \N__6494\,
            I => \N__6421\
        );

    \I__1368\ : ClkMux
    port map (
            O => \N__6493\,
            I => \N__6421\
        );

    \I__1367\ : ClkMux
    port map (
            O => \N__6492\,
            I => \N__6421\
        );

    \I__1366\ : ClkMux
    port map (
            O => \N__6491\,
            I => \N__6421\
        );

    \I__1365\ : ClkMux
    port map (
            O => \N__6490\,
            I => \N__6421\
        );

    \I__1364\ : ClkMux
    port map (
            O => \N__6489\,
            I => \N__6421\
        );

    \I__1363\ : ClkMux
    port map (
            O => \N__6488\,
            I => \N__6421\
        );

    \I__1362\ : ClkMux
    port map (
            O => \N__6487\,
            I => \N__6421\
        );

    \I__1361\ : ClkMux
    port map (
            O => \N__6486\,
            I => \N__6421\
        );

    \I__1360\ : ClkMux
    port map (
            O => \N__6485\,
            I => \N__6421\
        );

    \I__1359\ : ClkMux
    port map (
            O => \N__6484\,
            I => \N__6421\
        );

    \I__1358\ : GlobalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1357\ : gio2CtrlBuf
    port map (
            O => \N__6418\,
            I => \i_Clk_c_g\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6411\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6408\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6411\,
            I => \r_count_1hzZ0Z_14\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6408\,
            I => \r_count_1hzZ0Z_14\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6399\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6396\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6399\,
            I => \r_count_1hzZ0Z_22\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6396\,
            I => \r_count_1hzZ0Z_22\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__6391\,
            I => \N__6387\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6384\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6381\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6384\,
            I => \r_count_1hzZ0Z_9\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6381\,
            I => \r_count_1hzZ0Z_9\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6376\,
            I => \N__6372\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6375\,
            I => \N__6369\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__6372\,
            I => \r_count_1hzZ0Z_16\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6369\,
            I => \r_count_1hzZ0Z_16\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__6355\,
            I => \o_LED_43_5_and\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6348\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6345\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6348\,
            I => \r_count_1hzZ0Z_25\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6345\,
            I => \r_count_1hzZ0Z_25\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6340\,
            I => \N__6336\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6333\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6336\,
            I => \r_count_1hzZ0Z_26\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6333\,
            I => \r_count_1hzZ0Z_26\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__6328\,
            I => \N__6324\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6321\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6318\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6321\,
            I => \r_count_1hzZ0Z_24\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6318\,
            I => \r_count_1hzZ0Z_24\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6309\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6306\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6309\,
            I => \r_count_1hzZ0Z_27\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6306\,
            I => \r_count_1hzZ0Z_27\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6295\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1315\ : Span4Mux_v
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__6289\,
            I => \o_LED_43_6_and\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6282\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6279\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6274\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6274\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__6274\,
            I => \r_count_10hzZ0Z_19\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6271\,
            I => un2_r_count_10hz_1_cry_18
        );

    \I__1307\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6264\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6260\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6264\,
            I => \N__6257\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6254\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6260\,
            I => \r_count_10hzZ0Z_20\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__6257\,
            I => \r_count_10hzZ0Z_20\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6254\,
            I => \r_count_10hzZ0Z_20\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6244\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6244\,
            I => \N__6241\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__6241\,
            I => \un2_r_count_10hz_1_cry_19_THRU_CO\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6238\,
            I => un2_r_count_10hz_1_cry_19
        );

    \I__1296\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6231\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6228\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6231\,
            I => \N__6225\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6228\,
            I => \r_count_10hzZ0Z_21\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__6225\,
            I => \r_count_10hzZ0Z_21\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6220\,
            I => un2_r_count_10hz_1_cry_20
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6210\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6207\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6210\,
            I => \N__6204\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6207\,
            I => \r_count_10hzZ0Z_22\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__6204\,
            I => \r_count_10hzZ0Z_22\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6199\,
            I => un2_r_count_10hz_1_cry_21
        );

    \I__1283\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6192\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6189\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6192\,
            I => \r_count_10hzZ0Z_23\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6189\,
            I => \r_count_10hzZ0Z_23\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6184\,
            I => un2_r_count_10hz_1_cry_22
        );

    \I__1278\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6177\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6174\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6177\,
            I => \r_count_10hzZ0Z_24\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6174\,
            I => \r_count_10hzZ0Z_24\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6169\,
            I => un2_r_count_10hz_1_cry_23
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6166\,
            I => \N__6162\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6159\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6156\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6159\,
            I => \r_count_10hzZ0Z_25\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__6156\,
            I => \r_count_10hzZ0Z_25\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6151\,
            I => \bfn_12_6_0_\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6144\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6141\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6144\,
            I => \r_count_10hzZ0Z_26\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6141\,
            I => \r_count_10hzZ0Z_26\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6136\,
            I => un2_r_count_10hz_1_cry_25
        );

    \I__1262\ : InMux
    port map (
            O => \N__6133\,
            I => un2_r_count_10hz_1_cry_9
        );

    \I__1261\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6126\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6123\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6126\,
            I => \N__6120\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6123\,
            I => \r_count_10hzZ0Z_11\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__6120\,
            I => \r_count_10hzZ0Z_11\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6115\,
            I => un2_r_count_10hz_1_cry_10
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__6112\,
            I => \N__6107\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6104\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6101\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6098\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6104\,
            I => \r_count_10hzZ0Z_12\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6101\,
            I => \r_count_10hzZ0Z_12\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6098\,
            I => \r_count_10hzZ0Z_12\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6088\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6088\,
            I => \un2_r_count_10hz_1_cry_11_THRU_CO\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6085\,
            I => un2_r_count_10hz_1_cry_11
        );

    \I__1245\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6078\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6075\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6078\,
            I => \r_count_10hzZ0Z_13\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6075\,
            I => \r_count_10hzZ0Z_13\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6070\,
            I => un2_r_count_10hz_1_cry_12
        );

    \I__1240\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6063\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6060\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6063\,
            I => \r_count_10hzZ0Z_14\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6060\,
            I => \r_count_10hzZ0Z_14\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6055\,
            I => un2_r_count_10hz_1_cry_13
        );

    \I__1235\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6048\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6045\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6048\,
            I => \r_count_10hzZ0Z_15\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6045\,
            I => \r_count_10hzZ0Z_15\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6040\,
            I => un2_r_count_10hz_1_cry_14
        );

    \I__1230\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6032\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6029\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6026\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6032\,
            I => \r_count_10hzZ0Z_16\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6029\,
            I => \r_count_10hzZ0Z_16\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6026\,
            I => \r_count_10hzZ0Z_16\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6016\,
            I => \un2_r_count_10hz_1_cry_15_THRU_CO\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6013\,
            I => un2_r_count_10hz_1_cry_15
        );

    \I__1221\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6006\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6002\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6006\,
            I => \N__5999\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5996\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6002\,
            I => \r_count_10hzZ0Z_17\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__5999\,
            I => \r_count_10hzZ0Z_17\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5996\,
            I => \r_count_10hzZ0Z_17\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5986\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5986\,
            I => \N__5983\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__5983\,
            I => \un2_r_count_10hz_1_cry_16_THRU_CO\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5980\,
            I => \bfn_12_5_0_\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5973\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5970\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5967\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5970\,
            I => \r_count_10hzZ0Z_18\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5967\,
            I => \r_count_10hzZ0Z_18\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5962\,
            I => un2_r_count_10hz_1_cry_17
        );

    \I__1204\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5955\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5952\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5955\,
            I => \r_count_10hzZ0Z_2\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5952\,
            I => \r_count_10hzZ0Z_2\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5947\,
            I => un2_r_count_10hz_1_cry_1
        );

    \I__1199\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5940\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5937\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5940\,
            I => \r_count_10hzZ0Z_3\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5937\,
            I => \r_count_10hzZ0Z_3\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5932\,
            I => un2_r_count_10hz_1_cry_2
        );

    \I__1194\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5924\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5921\
        );

    \I__1192\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5918\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5924\,
            I => \r_count_10hzZ0Z_4\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5921\,
            I => \r_count_10hzZ0Z_4\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5918\,
            I => \r_count_10hzZ0Z_4\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5908\,
            I => \un2_r_count_10hz_1_cry_3_THRU_CO\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5905\,
            I => un2_r_count_10hz_1_cry_3
        );

    \I__1185\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5898\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5895\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5898\,
            I => \r_count_10hzZ0Z_5\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5895\,
            I => \r_count_10hzZ0Z_5\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5890\,
            I => un2_r_count_10hz_1_cry_4
        );

    \I__1180\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5882\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5879\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5876\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5882\,
            I => \r_count_10hzZ0Z_6\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5879\,
            I => \r_count_10hzZ0Z_6\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5876\,
            I => \r_count_10hzZ0Z_6\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5866\,
            I => \un2_r_count_10hz_1_cry_5_THRU_CO\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5863\,
            I => un2_r_count_10hz_1_cry_5
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__5860\,
            I => \N__5856\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5850\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5850\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5847\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5850\,
            I => \r_count_10hzZ0Z_7\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5847\,
            I => \r_count_10hzZ0Z_7\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5839\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5839\,
            I => \un2_r_count_10hz_1_cry_6_THRU_CO\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5836\,
            I => un2_r_count_10hz_1_cry_6
        );

    \I__1162\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5829\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5826\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5829\,
            I => \r_count_10hzZ0Z_8\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5826\,
            I => \r_count_10hzZ0Z_8\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5821\,
            I => un2_r_count_10hz_1_cry_7
        );

    \I__1157\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5813\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5810\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5807\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5813\,
            I => \r_count_10hzZ0Z_9\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5810\,
            I => \r_count_10hzZ0Z_9\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5807\,
            I => \r_count_10hzZ0Z_9\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5797\,
            I => \un2_r_count_10hz_1_cry_8_THRU_CO\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5794\,
            I => \bfn_12_4_0_\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__5791\,
            I => \N__5788\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5784\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5781\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5778\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5781\,
            I => \r_count_10hzZ0Z_10\
        );

    \I__1143\ : Odrv12
    port map (
            O => \N__5778\,
            I => \r_count_10hzZ0Z_10\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5767\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5767\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5767\,
            I => \r_count_1hzZ0Z_31\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__5764\,
            I => \N__5760\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__5763\,
            I => \N__5757\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5752\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5752\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5752\,
            I => \r_count_1hzZ0Z_28\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5743\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5743\,
            I => \r_count_1hzZ0Z_30\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__1128\ : Span4Mux_h
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__5728\,
            I => \o_LED_43_7_and\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__5725\,
            I => \N__5717\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__5724\,
            I => \N__5711\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__5723\,
            I => \N__5708\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5722\,
            I => \N__5705\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__5721\,
            I => \N__5702\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5695\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5695\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5695\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5715\,
            I => \N__5682\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5682\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5682\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5708\,
            I => \N__5682\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5682\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5682\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5695\,
            I => \o_LED_13_THRU_CO\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5682\,
            I => \o_LED_13_THRU_CO\
        );

    \I__1110\ : CascadeMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5671\,
            I => \o_LED_13_0_and\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5662\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5662\,
            I => \o_LED_13_3_and\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5656\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5656\,
            I => \o_LED_13_2_and\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__5653\,
            I => \N__5649\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__5652\,
            I => \N__5645\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5637\
        );

    \I__1099\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5637\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5637\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5634\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5637\,
            I => \r_count_10hzZ0Z_0\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5634\,
            I => \r_count_10hzZ0Z_0\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5622\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5622\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__5627\,
            I => \N__5619\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5616\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5613\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__5616\,
            I => \r_count_10hzZ0Z_1\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5613\,
            I => \r_count_10hzZ0Z_1\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5608\,
            I => un2_r_count_1hz_1_cry_22
        );

    \I__1086\ : InMux
    port map (
            O => \N__5605\,
            I => un2_r_count_1hz_1_cry_23
        );

    \I__1085\ : InMux
    port map (
            O => \N__5602\,
            I => \bfn_11_12_0_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5599\,
            I => un2_r_count_1hz_1_cry_25
        );

    \I__1083\ : InMux
    port map (
            O => \N__5596\,
            I => un2_r_count_1hz_1_cry_26
        );

    \I__1082\ : InMux
    port map (
            O => \N__5593\,
            I => un2_r_count_1hz_1_cry_27
        );

    \I__1081\ : InMux
    port map (
            O => \N__5590\,
            I => un2_r_count_1hz_1_cry_28
        );

    \I__1080\ : InMux
    port map (
            O => \N__5587\,
            I => un2_r_count_1hz_1_cry_29
        );

    \I__1079\ : InMux
    port map (
            O => \N__5584\,
            I => un2_r_count_1hz_1_cry_30
        );

    \I__1078\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5575\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5575\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5575\,
            I => \r_count_1hzZ0Z_29\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__5566\,
            I => \un2_r_count_1hz_1_cry_14_THRU_CO\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5563\,
            I => un2_r_count_1hz_1_cry_14
        );

    \I__1071\ : InMux
    port map (
            O => \N__5560\,
            I => un2_r_count_1hz_1_cry_15
        );

    \I__1070\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5552\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__5556\,
            I => \N__5549\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5546\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5543\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5540\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5546\,
            I => \r_count_1hzZ0Z_17\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5543\,
            I => \r_count_1hzZ0Z_17\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5540\,
            I => \r_count_1hzZ0Z_17\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__5524\,
            I => \un2_r_count_1hz_1_cry_16_THRU_CO\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5521\,
            I => \bfn_11_11_0_\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5514\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5511\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5514\,
            I => \N__5505\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5505\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5502\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__5505\,
            I => \r_count_1hzZ0Z_18\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5502\,
            I => \r_count_1hzZ0Z_18\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__1048\ : Span4Mux_h
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__5488\,
            I => \un2_r_count_1hz_1_cry_17_THRU_CO\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5485\,
            I => un2_r_count_1hz_1_cry_17
        );

    \I__1045\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5478\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5474\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5478\,
            I => \N__5471\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5468\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5474\,
            I => \r_count_1hzZ0Z_19\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__5471\,
            I => \r_count_1hzZ0Z_19\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5468\,
            I => \r_count_1hzZ0Z_19\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__1036\ : Span4Mux_h
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__5452\,
            I => \un2_r_count_1hz_1_cry_18_THRU_CO\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5449\,
            I => un2_r_count_1hz_1_cry_18
        );

    \I__1033\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5442\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5438\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5435\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5432\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5438\,
            I => \r_count_1hzZ0Z_20\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__5435\,
            I => \r_count_1hzZ0Z_20\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5432\,
            I => \r_count_1hzZ0Z_20\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5422\,
            I => \N__5419\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__5419\,
            I => \un2_r_count_1hz_1_cry_19_THRU_CO\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5416\,
            I => un2_r_count_1hz_1_cry_19
        );

    \I__1022\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5408\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__5412\,
            I => \N__5405\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5402\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5399\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5396\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5402\,
            I => \r_count_1hzZ0Z_21\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__5399\,
            I => \r_count_1hzZ0Z_21\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5396\,
            I => \r_count_1hzZ0Z_21\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1012\ : Odrv4
    port map (
            O => \N__5383\,
            I => \un2_r_count_1hz_1_cry_20_THRU_CO\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5380\,
            I => un2_r_count_1hz_1_cry_20
        );

    \I__1010\ : InMux
    port map (
            O => \N__5377\,
            I => un2_r_count_1hz_1_cry_21
        );

    \I__1009\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5369\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5366\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5363\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5369\,
            I => \N__5360\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5357\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5363\,
            I => \r_count_1hzZ0Z_23\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__5360\,
            I => \r_count_1hzZ0Z_23\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__5357\,
            I => \r_count_1hzZ0Z_23\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__5344\,
            I => \un2_r_count_1hz_1_cry_22_THRU_CO\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__5341\,
            I => \N__5338\
        );

    \I__997\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5334\
        );

    \I__996\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5331\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5334\,
            I => \r_count_1hzZ0Z_7\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5331\,
            I => \r_count_1hzZ0Z_7\
        );

    \I__993\ : InMux
    port map (
            O => \N__5326\,
            I => un2_r_count_1hz_1_cry_6
        );

    \I__992\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5319\
        );

    \I__991\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5316\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5319\,
            I => \r_count_1hzZ0Z_8\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5316\,
            I => \r_count_1hzZ0Z_8\
        );

    \I__988\ : InMux
    port map (
            O => \N__5311\,
            I => un2_r_count_1hz_1_cry_7
        );

    \I__987\ : InMux
    port map (
            O => \N__5308\,
            I => \bfn_11_10_0_\
        );

    \I__986\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5300\
        );

    \I__985\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5297\
        );

    \I__984\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5294\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5289\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5289\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5294\,
            I => \r_count_1hzZ0Z_10\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__5289\,
            I => \r_count_1hzZ0Z_10\
        );

    \I__979\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5281\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__977\ : Span4Mux_h
    port map (
            O => \N__5278\,
            I => \N__5275\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__5275\,
            I => \un2_r_count_1hz_1_cry_9_THRU_CO\
        );

    \I__975\ : InMux
    port map (
            O => \N__5272\,
            I => un2_r_count_1hz_1_cry_9
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__5269\,
            I => \N__5264\
        );

    \I__973\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5261\
        );

    \I__972\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5258\
        );

    \I__971\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5255\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5261\,
            I => \N__5252\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5258\,
            I => \r_count_1hzZ0Z_11\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5255\,
            I => \r_count_1hzZ0Z_11\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__5252\,
            I => \r_count_1hzZ0Z_11\
        );

    \I__966\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__964\ : Span4Mux_h
    port map (
            O => \N__5239\,
            I => \N__5236\
        );

    \I__963\ : Odrv4
    port map (
            O => \N__5236\,
            I => \un2_r_count_1hz_1_cry_10_THRU_CO\
        );

    \I__962\ : InMux
    port map (
            O => \N__5233\,
            I => un2_r_count_1hz_1_cry_10
        );

    \I__961\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5226\
        );

    \I__960\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5222\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5219\
        );

    \I__958\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5216\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5222\,
            I => \r_count_1hzZ0Z_12\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__5219\,
            I => \r_count_1hzZ0Z_12\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5216\,
            I => \r_count_1hzZ0Z_12\
        );

    \I__954\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5206\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__5200\,
            I => \un2_r_count_1hz_1_cry_11_THRU_CO\
        );

    \I__950\ : InMux
    port map (
            O => \N__5197\,
            I => un2_r_count_1hz_1_cry_11
        );

    \I__949\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5189\
        );

    \I__948\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5184\
        );

    \I__947\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5184\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5189\,
            I => \N__5181\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5184\,
            I => \r_count_1hzZ0Z_13\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__5181\,
            I => \r_count_1hzZ0Z_13\
        );

    \I__943\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__5170\,
            I => \un2_r_count_1hz_1_cry_12_THRU_CO\
        );

    \I__940\ : InMux
    port map (
            O => \N__5167\,
            I => un2_r_count_1hz_1_cry_12
        );

    \I__939\ : InMux
    port map (
            O => \N__5164\,
            I => un2_r_count_1hz_1_cry_13
        );

    \I__938\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5154\
        );

    \I__937\ : InMux
    port map (
            O => \N__5160\,
            I => \N__5154\
        );

    \I__936\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5151\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5146\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5146\,
            I => \r_count_1hzZ0Z_15\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__931\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5137\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__929\ : Span4Mux_h
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__5131\,
            I => \o_LED_43_4_and\
        );

    \I__927\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5124\
        );

    \I__926\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5121\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5124\,
            I => \N__5117\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5121\,
            I => \N__5113\
        );

    \I__923\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5110\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__5117\,
            I => \N__5107\
        );

    \I__921\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5104\
        );

    \I__920\ : Span4Mux_s3_h
    port map (
            O => \N__5113\,
            I => \N__5101\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5110\,
            I => \r_count_1hzZ0Z_0\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__5107\,
            I => \r_count_1hzZ0Z_0\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5104\,
            I => \r_count_1hzZ0Z_0\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__5101\,
            I => \r_count_1hzZ0Z_0\
        );

    \I__915\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5089\,
            I => \N__5084\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \N__5081\
        );

    \I__912\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5078\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__5084\,
            I => \N__5075\
        );

    \I__910\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5072\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5078\,
            I => \r_count_1hzZ0Z_1\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__5075\,
            I => \r_count_1hzZ0Z_1\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5072\,
            I => \r_count_1hzZ0Z_1\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__5065\,
            I => \N__5062\
        );

    \I__905\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5059\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__903\ : Span4Mux_h
    port map (
            O => \N__5056\,
            I => \N__5052\
        );

    \I__902\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__5052\,
            I => \r_count_1hzZ0Z_2\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5049\,
            I => \r_count_1hzZ0Z_2\
        );

    \I__899\ : InMux
    port map (
            O => \N__5044\,
            I => un2_r_count_1hz_1_cry_1
        );

    \I__898\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5034\
        );

    \I__896\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5031\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__5034\,
            I => \N__5028\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5031\,
            I => \r_count_1hzZ0Z_3\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__5028\,
            I => \r_count_1hzZ0Z_3\
        );

    \I__892\ : InMux
    port map (
            O => \N__5023\,
            I => un2_r_count_1hz_1_cry_2
        );

    \I__891\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5016\
        );

    \I__890\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5016\,
            I => \r_count_1hzZ0Z_4\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5013\,
            I => \r_count_1hzZ0Z_4\
        );

    \I__887\ : InMux
    port map (
            O => \N__5008\,
            I => un2_r_count_1hz_1_cry_3
        );

    \I__886\ : InMux
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5002\,
            I => \N__4997\
        );

    \I__884\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4992\
        );

    \I__883\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4992\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__4997\,
            I => \N__4989\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4992\,
            I => \r_count_1hzZ0Z_5\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4989\,
            I => \r_count_1hzZ0Z_5\
        );

    \I__879\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__877\ : Span4Mux_v
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__876\ : Odrv4
    port map (
            O => \N__4975\,
            I => \un2_r_count_1hz_1_cry_4_THRU_CO\
        );

    \I__875\ : InMux
    port map (
            O => \N__4972\,
            I => un2_r_count_1hz_1_cry_4
        );

    \I__874\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4965\
        );

    \I__873\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4962\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4965\,
            I => \r_count_1hzZ0Z_6\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4962\,
            I => \r_count_1hzZ0Z_6\
        );

    \I__870\ : InMux
    port map (
            O => \N__4957\,
            I => un2_r_count_1hz_1_cry_5
        );

    \I__869\ : IoInMux
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__867\ : Span4Mux_s1_h
    port map (
            O => \N__4948\,
            I => \N__4944\
        );

    \I__866\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4941\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4944\,
            I => \o_LED_1_c\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4941\,
            I => \o_LED_1_c\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__862\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__860\ : Odrv12
    port map (
            O => \N__4927\,
            I => \o_LED_13_4_and\
        );

    \I__859\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__4918\,
            I => \o_LED_13_5_and\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__855\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__853\ : Odrv12
    port map (
            O => \N__4906\,
            I => \o_LED_13_6_and\
        );

    \I__852\ : CascadeMux
    port map (
            O => \N__4903\,
            I => \N__4900\
        );

    \I__851\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__849\ : Odrv12
    port map (
            O => \N__4894\,
            I => \o_LED_13_7_and\
        );

    \I__848\ : InMux
    port map (
            O => \N__4891\,
            I => \bfn_11_2_0_\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__4888\,
            I => \o_LED_13_THRU_CO_cascade_\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4885\,
            I => \N__4882\
        );

    \I__845\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4879\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4879\,
            I => \o_LED_13_1_and\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__4876\,
            I => \N__4869\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__4875\,
            I => \N__4864\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \N__4860\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \N__4855\
        );

    \I__839\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4849\
        );

    \I__838\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4844\
        );

    \I__837\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4844\
        );

    \I__836\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4831\
        );

    \I__835\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4831\
        );

    \I__834\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4831\
        );

    \I__833\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4831\
        );

    \I__832\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4831\
        );

    \I__831\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4831\
        );

    \I__830\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4822\
        );

    \I__829\ : InMux
    port map (
            O => \N__4854\,
            I => \N__4822\
        );

    \I__828\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4822\
        );

    \I__827\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4822\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4849\,
            I => \o_LED_43_THRU_CO\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4844\,
            I => \o_LED_43_THRU_CO\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4831\,
            I => \o_LED_43_THRU_CO\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4822\,
            I => \o_LED_43_THRU_CO\
        );

    \I__822\ : InMux
    port map (
            O => \N__4813\,
            I => \bfn_9_10_0_\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \o_LED_43_THRU_CO_cascade_\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__819\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4801\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4801\,
            I => \o_LED_43_1_and\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__816\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4792\,
            I => \o_LED_43_2_and\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__813\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4782\
        );

    \I__812\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4779\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4779\,
            I => \r_count_5hzZ0Z_28\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__4776\,
            I => \r_count_5hzZ0Z_28\
        );

    \I__808\ : InMux
    port map (
            O => \N__4771\,
            I => un2_r_count_5hz_1_cry_27
        );

    \I__807\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4764\
        );

    \I__806\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4764\,
            I => \r_count_5hzZ0Z_29\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4761\,
            I => \r_count_5hzZ0Z_29\
        );

    \I__803\ : InMux
    port map (
            O => \N__4756\,
            I => un2_r_count_5hz_1_cry_28
        );

    \I__802\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4749\
        );

    \I__801\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4749\,
            I => \r_count_5hzZ0Z_30\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4746\,
            I => \r_count_5hzZ0Z_30\
        );

    \I__798\ : InMux
    port map (
            O => \N__4741\,
            I => un2_r_count_5hz_1_cry_29
        );

    \I__797\ : InMux
    port map (
            O => \N__4738\,
            I => un2_r_count_5hz_1_cry_30
        );

    \I__796\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4731\
        );

    \I__795\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4731\,
            I => \r_count_5hzZ0Z_31\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4728\,
            I => \r_count_5hzZ0Z_31\
        );

    \I__792\ : CascadeMux
    port map (
            O => \N__4723\,
            I => \N__4720\
        );

    \I__791\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4717\,
            I => \o_LED_43_0_and\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4714\,
            I => \N__4711\
        );

    \I__788\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4708\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4708\,
            I => \o_LED_43_3_and\
        );

    \I__786\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4701\
        );

    \I__785\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4698\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4701\,
            I => \r_count_5hzZ0Z_20\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4698\,
            I => \r_count_5hzZ0Z_20\
        );

    \I__782\ : InMux
    port map (
            O => \N__4693\,
            I => un2_r_count_5hz_1_cry_19
        );

    \I__781\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4686\
        );

    \I__780\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4683\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4686\,
            I => \N__4680\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4683\,
            I => \r_count_5hzZ0Z_21\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__4680\,
            I => \r_count_5hzZ0Z_21\
        );

    \I__776\ : InMux
    port map (
            O => \N__4675\,
            I => un2_r_count_5hz_1_cry_20
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__4672\,
            I => \N__4668\
        );

    \I__774\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4665\
        );

    \I__773\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4662\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4665\,
            I => \r_count_5hzZ0Z_22\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4662\,
            I => \r_count_5hzZ0Z_22\
        );

    \I__770\ : InMux
    port map (
            O => \N__4657\,
            I => un2_r_count_5hz_1_cry_21
        );

    \I__769\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4650\
        );

    \I__768\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4647\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4650\,
            I => \N__4642\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4647\,
            I => \N__4642\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__4642\,
            I => \r_count_5hzZ0Z_23\
        );

    \I__764\ : InMux
    port map (
            O => \N__4639\,
            I => un2_r_count_5hz_1_cry_22
        );

    \I__763\ : InMux
    port map (
            O => \N__4636\,
            I => \N__4632\
        );

    \I__762\ : InMux
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4632\,
            I => \r_count_5hzZ0Z_24\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4629\,
            I => \r_count_5hzZ0Z_24\
        );

    \I__759\ : InMux
    port map (
            O => \N__4624\,
            I => un2_r_count_5hz_1_cry_23
        );

    \I__758\ : InMux
    port map (
            O => \N__4621\,
            I => \N__4617\
        );

    \I__757\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4614\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__4617\,
            I => \r_count_5hzZ0Z_25\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4614\,
            I => \r_count_5hzZ0Z_25\
        );

    \I__754\ : InMux
    port map (
            O => \N__4609\,
            I => \bfn_9_5_0_\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__4606\,
            I => \N__4602\
        );

    \I__752\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4599\
        );

    \I__751\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4596\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4599\,
            I => \r_count_5hzZ0Z_26\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4596\,
            I => \r_count_5hzZ0Z_26\
        );

    \I__748\ : InMux
    port map (
            O => \N__4591\,
            I => un2_r_count_5hz_1_cry_25
        );

    \I__747\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4584\
        );

    \I__746\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4581\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4584\,
            I => \r_count_5hzZ0Z_27\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__4581\,
            I => \r_count_5hzZ0Z_27\
        );

    \I__743\ : InMux
    port map (
            O => \N__4576\,
            I => un2_r_count_5hz_1_cry_26
        );

    \I__742\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4568\
        );

    \I__741\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4563\
        );

    \I__740\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4563\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4568\,
            I => \r_count_5hzZ0Z_12\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4563\,
            I => \r_count_5hzZ0Z_12\
        );

    \I__737\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4555\,
            I => \un2_r_count_5hz_1_cry_11_THRU_CO\
        );

    \I__735\ : InMux
    port map (
            O => \N__4552\,
            I => un2_r_count_5hz_1_cry_11
        );

    \I__734\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4545\
        );

    \I__733\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4542\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4545\,
            I => \r_count_5hzZ0Z_13\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4542\,
            I => \r_count_5hzZ0Z_13\
        );

    \I__730\ : InMux
    port map (
            O => \N__4537\,
            I => un2_r_count_5hz_1_cry_12
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__4534\,
            I => \N__4529\
        );

    \I__728\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4526\
        );

    \I__727\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4523\
        );

    \I__726\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4520\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4526\,
            I => \r_count_5hzZ0Z_14\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__4523\,
            I => \r_count_5hzZ0Z_14\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4520\,
            I => \r_count_5hzZ0Z_14\
        );

    \I__722\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4510\,
            I => \un2_r_count_5hz_1_cry_13_THRU_CO\
        );

    \I__720\ : InMux
    port map (
            O => \N__4507\,
            I => un2_r_count_5hz_1_cry_13
        );

    \I__719\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4499\
        );

    \I__718\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4494\
        );

    \I__717\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4494\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4499\,
            I => \r_count_5hzZ0Z_15\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4494\,
            I => \r_count_5hzZ0Z_15\
        );

    \I__714\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4486\,
            I => \un2_r_count_5hz_1_cry_14_THRU_CO\
        );

    \I__712\ : InMux
    port map (
            O => \N__4483\,
            I => un2_r_count_5hz_1_cry_14
        );

    \I__711\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4475\
        );

    \I__710\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4472\
        );

    \I__709\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4469\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4466\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4472\,
            I => \r_count_5hzZ0Z_16\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4469\,
            I => \r_count_5hzZ0Z_16\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__4466\,
            I => \r_count_5hzZ0Z_16\
        );

    \I__704\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4456\,
            I => \un2_r_count_5hz_1_cry_15_THRU_CO\
        );

    \I__702\ : InMux
    port map (
            O => \N__4453\,
            I => un2_r_count_5hz_1_cry_15
        );

    \I__701\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4445\
        );

    \I__700\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4442\
        );

    \I__699\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4439\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4445\,
            I => \r_count_5hzZ0Z_17\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4442\,
            I => \r_count_5hzZ0Z_17\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4439\,
            I => \r_count_5hzZ0Z_17\
        );

    \I__695\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4429\,
            I => \un2_r_count_5hz_1_cry_16_THRU_CO\
        );

    \I__693\ : InMux
    port map (
            O => \N__4426\,
            I => \bfn_9_4_0_\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__4423\,
            I => \N__4419\
        );

    \I__691\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4416\
        );

    \I__690\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4408\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4408\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__4408\,
            I => \r_count_5hzZ0Z_18\
        );

    \I__686\ : InMux
    port map (
            O => \N__4405\,
            I => un2_r_count_5hz_1_cry_17
        );

    \I__685\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4398\
        );

    \I__684\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4395\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4398\,
            I => \r_count_5hzZ0Z_19\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4395\,
            I => \r_count_5hzZ0Z_19\
        );

    \I__681\ : InMux
    port map (
            O => \N__4390\,
            I => un2_r_count_5hz_1_cry_18
        );

    \I__680\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4380\
        );

    \I__679\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__678\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4377\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4380\,
            I => \r_count_5hzZ0Z_4\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4377\,
            I => \r_count_5hzZ0Z_4\
        );

    \I__675\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4369\,
            I => \un2_r_count_5hz_1_cry_3_THRU_CO\
        );

    \I__673\ : InMux
    port map (
            O => \N__4366\,
            I => un2_r_count_5hz_1_cry_3
        );

    \I__672\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4359\
        );

    \I__671\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4356\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4359\,
            I => \r_count_5hzZ0Z_5\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4356\,
            I => \r_count_5hzZ0Z_5\
        );

    \I__668\ : InMux
    port map (
            O => \N__4351\,
            I => un2_r_count_5hz_1_cry_4
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__666\ : InMux
    port map (
            O => \N__4345\,
            I => \N__4341\
        );

    \I__665\ : InMux
    port map (
            O => \N__4344\,
            I => \N__4338\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4341\,
            I => \r_count_5hzZ0Z_6\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4338\,
            I => \r_count_5hzZ0Z_6\
        );

    \I__662\ : InMux
    port map (
            O => \N__4333\,
            I => un2_r_count_5hz_1_cry_5
        );

    \I__661\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4325\
        );

    \I__660\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4322\
        );

    \I__659\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4319\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4325\,
            I => \r_count_5hzZ0Z_7\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4322\,
            I => \r_count_5hzZ0Z_7\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4319\,
            I => \r_count_5hzZ0Z_7\
        );

    \I__655\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4309\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4309\,
            I => \un2_r_count_5hz_1_cry_6_THRU_CO\
        );

    \I__653\ : InMux
    port map (
            O => \N__4306\,
            I => un2_r_count_5hz_1_cry_6
        );

    \I__652\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4299\
        );

    \I__651\ : InMux
    port map (
            O => \N__4302\,
            I => \N__4296\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4299\,
            I => \r_count_5hzZ0Z_8\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4296\,
            I => \r_count_5hzZ0Z_8\
        );

    \I__648\ : InMux
    port map (
            O => \N__4291\,
            I => un2_r_count_5hz_1_cry_7
        );

    \I__647\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4284\
        );

    \I__646\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4284\,
            I => \r_count_5hzZ0Z_9\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4281\,
            I => \r_count_5hzZ0Z_9\
        );

    \I__643\ : InMux
    port map (
            O => \N__4276\,
            I => \bfn_9_3_0_\
        );

    \I__642\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4269\
        );

    \I__641\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4269\,
            I => \r_count_5hzZ0Z_10\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4266\,
            I => \r_count_5hzZ0Z_10\
        );

    \I__638\ : InMux
    port map (
            O => \N__4261\,
            I => un2_r_count_5hz_1_cry_9
        );

    \I__637\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4254\
        );

    \I__636\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4251\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4254\,
            I => \r_count_5hzZ0Z_11\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4251\,
            I => \r_count_5hzZ0Z_11\
        );

    \I__633\ : InMux
    port map (
            O => \N__4246\,
            I => un2_r_count_5hz_1_cry_10
        );

    \I__632\ : InMux
    port map (
            O => \N__4243\,
            I => un2_r_count_2hz_1_cry_30
        );

    \I__631\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4236\
        );

    \I__630\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4233\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4236\,
            I => \r_count_2hzZ0Z_31\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4233\,
            I => \r_count_2hzZ0Z_31\
        );

    \I__627\ : IoInMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N__4222\
        );

    \I__625\ : Span4Mux_s3_h
    port map (
            O => \N__4222\,
            I => \N__4218\
        );

    \I__624\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__4218\,
            I => \o_LED_4_c\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4215\,
            I => \o_LED_4_c\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__4210\,
            I => \N__4205\
        );

    \I__620\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4201\
        );

    \I__619\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4196\
        );

    \I__618\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4196\
        );

    \I__617\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4193\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4201\,
            I => \r_count_5hzZ0Z_0\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4196\,
            I => \r_count_5hzZ0Z_0\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4193\,
            I => \r_count_5hzZ0Z_0\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__4186\,
            I => \N__4181\
        );

    \I__612\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4176\
        );

    \I__611\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4176\
        );

    \I__610\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4173\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4176\,
            I => \r_count_5hzZ0Z_1\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4173\,
            I => \r_count_5hzZ0Z_1\
        );

    \I__607\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4161\
        );

    \I__605\ : InMux
    port map (
            O => \N__4164\,
            I => \N__4158\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__4161\,
            I => \r_count_5hzZ0Z_2\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4158\,
            I => \r_count_5hzZ0Z_2\
        );

    \I__602\ : InMux
    port map (
            O => \N__4153\,
            I => un2_r_count_5hz_1_cry_1
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__600\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4143\
        );

    \I__599\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4140\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4143\,
            I => \r_count_5hzZ0Z_3\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4140\,
            I => \r_count_5hzZ0Z_3\
        );

    \I__596\ : InMux
    port map (
            O => \N__4135\,
            I => un2_r_count_5hz_1_cry_2
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__4132\,
            I => \N__4127\
        );

    \I__594\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4124\
        );

    \I__593\ : InMux
    port map (
            O => \N__4130\,
            I => \N__4121\
        );

    \I__592\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4118\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4124\,
            I => \r_count_2hzZ0Z_22\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4121\,
            I => \r_count_2hzZ0Z_22\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4118\,
            I => \r_count_2hzZ0Z_22\
        );

    \I__588\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4108\,
            I => \un2_r_count_2hz_1_cry_21_THRU_CO\
        );

    \I__586\ : InMux
    port map (
            O => \N__4105\,
            I => un2_r_count_2hz_1_cry_21
        );

    \I__585\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4098\
        );

    \I__584\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4095\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4098\,
            I => \r_count_2hzZ0Z_23\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4095\,
            I => \r_count_2hzZ0Z_23\
        );

    \I__581\ : InMux
    port map (
            O => \N__4090\,
            I => un2_r_count_2hz_1_cry_22
        );

    \I__580\ : CascadeMux
    port map (
            O => \N__4087\,
            I => \N__4083\
        );

    \I__579\ : InMux
    port map (
            O => \N__4086\,
            I => \N__4080\
        );

    \I__578\ : InMux
    port map (
            O => \N__4083\,
            I => \N__4077\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4080\,
            I => \r_count_2hzZ0Z_24\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4077\,
            I => \r_count_2hzZ0Z_24\
        );

    \I__575\ : InMux
    port map (
            O => \N__4072\,
            I => un2_r_count_2hz_1_cry_23
        );

    \I__574\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4065\
        );

    \I__573\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4062\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4065\,
            I => \r_count_2hzZ0Z_25\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4062\,
            I => \r_count_2hzZ0Z_25\
        );

    \I__570\ : InMux
    port map (
            O => \N__4057\,
            I => \bfn_8_9_0_\
        );

    \I__569\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4050\
        );

    \I__568\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4047\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4050\,
            I => \N__4044\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4047\,
            I => \r_count_2hzZ0Z_26\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__4044\,
            I => \r_count_2hzZ0Z_26\
        );

    \I__564\ : InMux
    port map (
            O => \N__4039\,
            I => un2_r_count_2hz_1_cry_25
        );

    \I__563\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4032\
        );

    \I__562\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4029\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4032\,
            I => \r_count_2hzZ0Z_27\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4029\,
            I => \r_count_2hzZ0Z_27\
        );

    \I__559\ : InMux
    port map (
            O => \N__4024\,
            I => un2_r_count_2hz_1_cry_26
        );

    \I__558\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4017\
        );

    \I__557\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4014\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4017\,
            I => \r_count_2hzZ0Z_28\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4014\,
            I => \r_count_2hzZ0Z_28\
        );

    \I__554\ : InMux
    port map (
            O => \N__4009\,
            I => un2_r_count_2hz_1_cry_27
        );

    \I__553\ : InMux
    port map (
            O => \N__4006\,
            I => \N__4002\
        );

    \I__552\ : InMux
    port map (
            O => \N__4005\,
            I => \N__3999\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4002\,
            I => \r_count_2hzZ0Z_29\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3999\,
            I => \r_count_2hzZ0Z_29\
        );

    \I__549\ : InMux
    port map (
            O => \N__3994\,
            I => un2_r_count_2hz_1_cry_28
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3991\,
            I => \N__3987\
        );

    \I__547\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3984\
        );

    \I__546\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3981\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3984\,
            I => \r_count_2hzZ0Z_30\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3981\,
            I => \r_count_2hzZ0Z_30\
        );

    \I__543\ : InMux
    port map (
            O => \N__3976\,
            I => un2_r_count_2hz_1_cry_29
        );

    \I__542\ : InMux
    port map (
            O => \N__3973\,
            I => \N__3970\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3970\,
            I => \N__3965\
        );

    \I__540\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3962\
        );

    \I__539\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3959\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__3965\,
            I => \r_count_2hzZ0Z_14\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3962\,
            I => \r_count_2hzZ0Z_14\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3959\,
            I => \r_count_2hzZ0Z_14\
        );

    \I__535\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3949\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3949\,
            I => \un2_r_count_2hz_1_cry_13_THRU_CO\
        );

    \I__533\ : InMux
    port map (
            O => \N__3946\,
            I => un2_r_count_2hz_1_cry_13
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__3943\,
            I => \N__3939\
        );

    \I__531\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3936\
        );

    \I__530\ : InMux
    port map (
            O => \N__3939\,
            I => \N__3933\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3936\,
            I => \r_count_2hzZ0Z_15\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3933\,
            I => \r_count_2hzZ0Z_15\
        );

    \I__527\ : InMux
    port map (
            O => \N__3928\,
            I => un2_r_count_2hz_1_cry_14
        );

    \I__526\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3920\
        );

    \I__525\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3917\
        );

    \I__524\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3914\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3920\,
            I => \r_count_2hzZ0Z_16\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3917\,
            I => \r_count_2hzZ0Z_16\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3914\,
            I => \r_count_2hzZ0Z_16\
        );

    \I__520\ : InMux
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__3901\,
            I => \un2_r_count_2hz_1_cry_15_THRU_CO\
        );

    \I__517\ : InMux
    port map (
            O => \N__3898\,
            I => un2_r_count_2hz_1_cry_15
        );

    \I__516\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3892\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3892\,
            I => \N__3887\
        );

    \I__514\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3882\
        );

    \I__513\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3882\
        );

    \I__512\ : Odrv4
    port map (
            O => \N__3887\,
            I => \r_count_2hzZ0Z_17\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3882\,
            I => \r_count_2hzZ0Z_17\
        );

    \I__510\ : InMux
    port map (
            O => \N__3877\,
            I => \N__3874\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3874\,
            I => \N__3871\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__3871\,
            I => \un2_r_count_2hz_1_cry_16_THRU_CO\
        );

    \I__507\ : InMux
    port map (
            O => \N__3868\,
            I => \bfn_8_8_0_\
        );

    \I__506\ : InMux
    port map (
            O => \N__3865\,
            I => \N__3860\
        );

    \I__505\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3857\
        );

    \I__504\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3854\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3860\,
            I => \r_count_2hzZ0Z_18\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3857\,
            I => \r_count_2hzZ0Z_18\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3854\,
            I => \r_count_2hzZ0Z_18\
        );

    \I__500\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3844\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3844\,
            I => \un2_r_count_2hz_1_cry_17_THRU_CO\
        );

    \I__498\ : InMux
    port map (
            O => \N__3841\,
            I => un2_r_count_2hz_1_cry_17
        );

    \I__497\ : InMux
    port map (
            O => \N__3838\,
            I => \N__3833\
        );

    \I__496\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3830\
        );

    \I__495\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3827\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3833\,
            I => \r_count_2hzZ0Z_19\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3830\,
            I => \r_count_2hzZ0Z_19\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3827\,
            I => \r_count_2hzZ0Z_19\
        );

    \I__491\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3817\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3817\,
            I => \N__3814\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__3814\,
            I => \un2_r_count_2hz_1_cry_18_THRU_CO\
        );

    \I__488\ : InMux
    port map (
            O => \N__3811\,
            I => un2_r_count_2hz_1_cry_18
        );

    \I__487\ : InMux
    port map (
            O => \N__3808\,
            I => \N__3803\
        );

    \I__486\ : InMux
    port map (
            O => \N__3807\,
            I => \N__3800\
        );

    \I__485\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3797\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3803\,
            I => \r_count_2hzZ0Z_20\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3800\,
            I => \r_count_2hzZ0Z_20\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3797\,
            I => \r_count_2hzZ0Z_20\
        );

    \I__481\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3787\,
            I => \un2_r_count_2hz_1_cry_19_THRU_CO\
        );

    \I__479\ : InMux
    port map (
            O => \N__3784\,
            I => un2_r_count_2hz_1_cry_19
        );

    \I__478\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3777\
        );

    \I__477\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3774\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3777\,
            I => \r_count_2hzZ0Z_21\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3774\,
            I => \r_count_2hzZ0Z_21\
        );

    \I__474\ : InMux
    port map (
            O => \N__3769\,
            I => un2_r_count_2hz_1_cry_20
        );

    \I__473\ : InMux
    port map (
            O => \N__3766\,
            I => \N__3762\
        );

    \I__472\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3759\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3762\,
            I => \r_count_2hzZ0Z_6\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3759\,
            I => \r_count_2hzZ0Z_6\
        );

    \I__469\ : InMux
    port map (
            O => \N__3754\,
            I => un2_r_count_2hz_1_cry_5
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__467\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3744\
        );

    \I__466\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3741\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3744\,
            I => \r_count_2hzZ0Z_7\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3741\,
            I => \r_count_2hzZ0Z_7\
        );

    \I__463\ : InMux
    port map (
            O => \N__3736\,
            I => un2_r_count_2hz_1_cry_6
        );

    \I__462\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3729\
        );

    \I__461\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3726\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3729\,
            I => \r_count_2hzZ0Z_8\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3726\,
            I => \r_count_2hzZ0Z_8\
        );

    \I__458\ : InMux
    port map (
            O => \N__3721\,
            I => un2_r_count_2hz_1_cry_7
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__456\ : InMux
    port map (
            O => \N__3715\,
            I => \N__3708\
        );

    \I__455\ : InMux
    port map (
            O => \N__3714\,
            I => \N__3708\
        );

    \I__454\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3705\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3708\,
            I => \r_count_2hzZ0Z_9\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3705\,
            I => \r_count_2hzZ0Z_9\
        );

    \I__451\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3697\,
            I => \un2_r_count_2hz_1_cry_8_THRU_CO\
        );

    \I__449\ : InMux
    port map (
            O => \N__3694\,
            I => \bfn_8_7_0_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__3691\,
            I => \N__3687\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3690\,
            I => \N__3684\
        );

    \I__446\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3678\
        );

    \I__445\ : InMux
    port map (
            O => \N__3684\,
            I => \N__3678\
        );

    \I__444\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3675\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3678\,
            I => \N__3672\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3675\,
            I => \r_count_2hzZ0Z_10\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__3672\,
            I => \r_count_2hzZ0Z_10\
        );

    \I__440\ : InMux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3664\,
            I => \un2_r_count_2hz_1_cry_9_THRU_CO\
        );

    \I__438\ : InMux
    port map (
            O => \N__3661\,
            I => un2_r_count_2hz_1_cry_9
        );

    \I__437\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3653\
        );

    \I__436\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3648\
        );

    \I__435\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3648\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3653\,
            I => \r_count_2hzZ0Z_11\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__3648\,
            I => \r_count_2hzZ0Z_11\
        );

    \I__432\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3640\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3640\,
            I => \un2_r_count_2hz_1_cry_10_THRU_CO\
        );

    \I__430\ : InMux
    port map (
            O => \N__3637\,
            I => un2_r_count_2hz_1_cry_10
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__3634\,
            I => \N__3629\
        );

    \I__428\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3626\
        );

    \I__427\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3623\
        );

    \I__426\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3620\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3626\,
            I => \r_count_2hzZ0Z_12\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3623\,
            I => \r_count_2hzZ0Z_12\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3620\,
            I => \r_count_2hzZ0Z_12\
        );

    \I__422\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3610\,
            I => \un2_r_count_2hz_1_cry_11_THRU_CO\
        );

    \I__420\ : InMux
    port map (
            O => \N__3607\,
            I => un2_r_count_2hz_1_cry_11
        );

    \I__419\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3600\
        );

    \I__418\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3597\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3600\,
            I => \r_count_2hzZ0Z_13\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3597\,
            I => \r_count_2hzZ0Z_13\
        );

    \I__415\ : InMux
    port map (
            O => \N__3592\,
            I => un2_r_count_2hz_1_cry_12
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3589\,
            I => \N__3586\
        );

    \I__413\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3583\,
            I => \o_LED_23_6_and\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__410\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3574\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3574\,
            I => \o_LED_23_4_and\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3571\,
            I => \N__3564\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__3570\,
            I => \N__3560\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3569\,
            I => \N__3555\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3568\,
            I => \N__3551\
        );

    \I__404\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3538\
        );

    \I__403\ : InMux
    port map (
            O => \N__3564\,
            I => \N__3538\
        );

    \I__402\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3538\
        );

    \I__401\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3538\
        );

    \I__400\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3538\
        );

    \I__399\ : InMux
    port map (
            O => \N__3558\,
            I => \N__3538\
        );

    \I__398\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3531\
        );

    \I__397\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3531\
        );

    \I__396\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3531\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3538\,
            I => \o_LED_23_THRU_CO\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3531\,
            I => \o_LED_23_THRU_CO\
        );

    \I__393\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3520\
        );

    \I__392\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3515\
        );

    \I__391\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3515\
        );

    \I__390\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3512\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__3520\,
            I => \r_count_2hzZ0Z_0\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3515\,
            I => \r_count_2hzZ0Z_0\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3512\,
            I => \r_count_2hzZ0Z_0\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3505\,
            I => \N__3500\
        );

    \I__385\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3497\
        );

    \I__384\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3494\
        );

    \I__383\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3491\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3497\,
            I => \r_count_2hzZ0Z_1\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3494\,
            I => \r_count_2hzZ0Z_1\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3491\,
            I => \r_count_2hzZ0Z_1\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__3484\,
            I => \N__3480\
        );

    \I__378\ : InMux
    port map (
            O => \N__3483\,
            I => \N__3477\
        );

    \I__377\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3474\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3477\,
            I => \r_count_2hzZ0Z_2\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3474\,
            I => \r_count_2hzZ0Z_2\
        );

    \I__374\ : InMux
    port map (
            O => \N__3469\,
            I => un2_r_count_2hz_1_cry_1
        );

    \I__373\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3462\
        );

    \I__372\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3459\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__3462\,
            I => \r_count_2hzZ0Z_3\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3459\,
            I => \r_count_2hzZ0Z_3\
        );

    \I__369\ : InMux
    port map (
            O => \N__3454\,
            I => un2_r_count_2hz_1_cry_2
        );

    \I__368\ : InMux
    port map (
            O => \N__3451\,
            I => \N__3444\
        );

    \I__367\ : InMux
    port map (
            O => \N__3450\,
            I => \N__3444\
        );

    \I__366\ : InMux
    port map (
            O => \N__3449\,
            I => \N__3441\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3444\,
            I => \r_count_2hzZ0Z_4\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3441\,
            I => \r_count_2hzZ0Z_4\
        );

    \I__363\ : InMux
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3433\,
            I => \un2_r_count_2hz_1_cry_3_THRU_CO\
        );

    \I__361\ : InMux
    port map (
            O => \N__3430\,
            I => un2_r_count_2hz_1_cry_3
        );

    \I__360\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3423\
        );

    \I__359\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3420\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3423\,
            I => \r_count_2hzZ0Z_5\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3420\,
            I => \r_count_2hzZ0Z_5\
        );

    \I__356\ : InMux
    port map (
            O => \N__3415\,
            I => un2_r_count_2hz_1_cry_4
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \N__3409\
        );

    \I__354\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3406\,
            I => \o_LED_23_1_and\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \N__3400\
        );

    \I__351\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3397\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3397\,
            I => \o_LED_23_0_and\
        );

    \I__349\ : CascadeMux
    port map (
            O => \N__3394\,
            I => \N__3391\
        );

    \I__348\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3388\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3388\,
            I => \o_LED_23_7_and\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__3385\,
            I => \N__3382\
        );

    \I__345\ : InMux
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3379\,
            I => \o_LED_23_5_and\
        );

    \I__343\ : IoInMux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__341\ : Span4Mux_s3_h
    port map (
            O => \N__3370\,
            I => \N__3366\
        );

    \I__340\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3363\
        );

    \I__339\ : Odrv4
    port map (
            O => \N__3366\,
            I => \o_LED_2_c\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3363\,
            I => \o_LED_2_c\
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__3358\,
            I => \N__3349\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__3357\,
            I => \N__3345\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__3356\,
            I => \N__3342\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3355\,
            I => \N__3338\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__3354\,
            I => \N__3333\
        );

    \I__332\ : CascadeMux
    port map (
            O => \N__3353\,
            I => \N__3329\
        );

    \I__331\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3325\
        );

    \I__330\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3314\
        );

    \I__329\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3314\
        );

    \I__328\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3314\
        );

    \I__327\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3314\
        );

    \I__326\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3314\
        );

    \I__325\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3299\
        );

    \I__324\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3299\
        );

    \I__323\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3299\
        );

    \I__322\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3299\
        );

    \I__321\ : InMux
    port map (
            O => \N__3332\,
            I => \N__3299\
        );

    \I__320\ : InMux
    port map (
            O => \N__3329\,
            I => \N__3299\
        );

    \I__319\ : InMux
    port map (
            O => \N__3328\,
            I => \N__3299\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3325\,
            I => \o_LED_33_THRU_CO\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3314\,
            I => \o_LED_33_THRU_CO\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3299\,
            I => \o_LED_33_THRU_CO\
        );

    \I__315\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__314\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3286\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__3286\,
            I => \N__3283\
        );

    \I__312\ : Odrv4
    port map (
            O => \N__3283\,
            I => \o_LED_33_7_and\
        );

    \I__311\ : CascadeMux
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__310\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3274\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3274\,
            I => \o_LED_23_2_and\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__3271\,
            I => \N__3268\
        );

    \I__307\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__3265\,
            I => \o_LED_23_3_and\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__304\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3256\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3256\,
            I => \o_LED_33_5_and\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__3253\,
            I => \N__3250\
        );

    \I__301\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3247\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__3247\,
            I => \o_LED_33_0_and\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__298\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__3238\,
            I => \o_LED_33_6_and\
        );

    \I__296\ : InMux
    port map (
            O => \N__3235\,
            I => \bfn_7_4_0_\
        );

    \I__295\ : CascadeMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__294\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__3226\,
            I => \o_LED_33_4_and\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__291\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__3217\,
            I => \o_LED_33_3_and\
        );

    \I__289\ : InMux
    port map (
            O => \N__3214\,
            I => \bfn_6_8_0_\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__3211\,
            I => \o_LED_33_THRU_CO_cascade_\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__285\ : Span4Mux_s2_h
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__284\ : Span4Mux_h
    port map (
            O => \N__3199\,
            I => \N__3195\
        );

    \I__283\ : InMux
    port map (
            O => \N__3198\,
            I => \N__3192\
        );

    \I__282\ : Odrv4
    port map (
            O => \N__3195\,
            I => \o_LED_3_c\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__3192\,
            I => \o_LED_3_c\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__3187\,
            I => \N__3184\
        );

    \I__279\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3181\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__3181\,
            I => \o_LED_33_2_and\
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__3178\,
            I => \N__3175\
        );

    \I__276\ : InMux
    port map (
            O => \N__3175\,
            I => \N__3172\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__3172\,
            I => \o_LED_33_1_and\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_5hz_1_cry_8,
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_5hz_1_cry_16,
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_5hz_1_cry_24,
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_2hz_1_cry_8,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_2hz_1_cry_16,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_2hz_1_cry_24,
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_1hz_1_cry_8,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_1hz_1_cry_16,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_1hz_1_cry_24,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_3_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_10hz_1_cry_8,
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_10hz_1_cry_16,
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un2_r_count_10hz_1_cry_24,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \o_LED_43\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \o_LED_33\,
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \o_LED_23\,
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_11_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_1_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \o_LED_13\,
            carryinitout => \bfn_11_2_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \o_LED_33_0_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3253\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \o_LED_33_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_1_c_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3178\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_0\,
            carryout => \o_LED_33_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_2_c_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3187\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_1\,
            carryout => \o_LED_33_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_3_c_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3223\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_2\,
            carryout => \o_LED_33_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_4_c_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3232\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_3\,
            carryout => \o_LED_33_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_5_c_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3262\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_4\,
            carryout => \o_LED_33_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_6_c_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3244\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_5\,
            carryout => \o_LED_33_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_7_c_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3292\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_33_6\,
            carryout => \o_LED_33\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_THRU_LUT4_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3214\,
            lcout => \o_LED_33_THRU_CO\,
            ltout => \o_LED_33_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_17_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__3891\,
            in1 => \N__3877\,
            in2 => \N__3211\,
            in3 => \_gnd_net_\,
            lcout => \r_count_2hzZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LEDZ0Z_3_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3198\,
            in2 => \_gnd_net_\,
            in3 => \N__3352\,
            lcout => \o_LED_3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6484\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_2_c_RNO_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3863\,
            in1 => \N__3836\,
            in2 => \N__4132\,
            in3 => \N__3806\,
            lcout => \o_LED_33_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_1_c_RNO_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3890\,
            in1 => \N__3968\,
            in2 => \N__3634\,
            in3 => \N__3923\,
            lcout => \o_LED_33_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_0_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3403\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \o_LED_23_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_1_c_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_0\,
            carryout => \o_LED_23_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_2_c_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3280\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_1\,
            carryout => \o_LED_23_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_3_c_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3271\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_2\,
            carryout => \o_LED_23_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_4_c_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3580\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_3\,
            carryout => \o_LED_23_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_5_c_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_4\,
            carryout => \o_LED_23_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_6_c_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_5\,
            carryout => \o_LED_23_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_7_c_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3394\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_23_6\,
            carryout => \o_LED_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_THRU_LUT4_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3235\,
            lcout => \o_LED_23_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3526\,
            in2 => \_gnd_net_\,
            in3 => \N__3504\,
            lcout => \r_count_2hzZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_4_c_RNO_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3766\,
            in1 => \N__3427\,
            in2 => \N__3751\,
            in3 => \N__3732\,
            lcout => \o_LED_33_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_10_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__3667\,
            in1 => \_gnd_net_\,
            in2 => \N__3691\,
            in3 => \N__3341\,
            lcout => \r_count_2hzZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__3525\,
            in1 => \_gnd_net_\,
            in2 => \N__3358\,
            in3 => \_gnd_net_\,
            lcout => \r_count_2hzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_3_c_RNO_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3503\,
            in1 => \N__3524\,
            in2 => \N__3484\,
            in3 => \N__3465\,
            lcout => \o_LED_33_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_11_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3657\,
            in1 => \_gnd_net_\,
            in2 => \N__3356\,
            in3 => \N__3643\,
            lcout => \r_count_2hzZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_9_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__3700\,
            in1 => \_gnd_net_\,
            in2 => \N__3718\,
            in3 => \N__3348\,
            lcout => \r_count_2hzZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_5_c_RNO_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3604\,
            in1 => \N__4101\,
            in2 => \N__3943\,
            in3 => \N__3780\,
            lcout => \o_LED_33_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_0_c_RNO_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3714\,
            in1 => \N__3450\,
            in2 => \N__3690\,
            in3 => \N__3656\,
            lcout => \o_LED_33_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_4_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3451\,
            in1 => \_gnd_net_\,
            in2 => \N__3357\,
            in3 => \N__3436\,
            lcout => \r_count_2hzZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_16_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3907\,
            in1 => \N__3925\,
            in2 => \_gnd_net_\,
            in3 => \N__3332\,
            lcout => \r_count_2hzZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_14_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3952\,
            in1 => \_gnd_net_\,
            in2 => \N__3353\,
            in3 => \N__3973\,
            lcout => \r_count_2hzZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_19_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3820\,
            in1 => \N__3838\,
            in2 => \_gnd_net_\,
            in3 => \N__3336\,
            lcout => \r_count_2hzZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_6_c_RNO_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4054\,
            in1 => \N__4068\,
            in2 => \N__4087\,
            in3 => \N__4035\,
            lcout => \o_LED_33_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_20_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3790\,
            in1 => \N__3808\,
            in2 => \_gnd_net_\,
            in3 => \N__3337\,
            lcout => \r_count_2hzZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_18_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3847\,
            in1 => \_gnd_net_\,
            in2 => \N__3354\,
            in3 => \N__3865\,
            lcout => \r_count_2hzZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_12_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3613\,
            in1 => \N__3633\,
            in2 => \_gnd_net_\,
            in3 => \N__3328\,
            lcout => \r_count_2hzZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_22_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4111\,
            in2 => \N__3355\,
            in3 => \N__4131\,
            lcout => \r_count_2hzZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_33_7_c_RNO_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4020\,
            in1 => \N__4239\,
            in2 => \N__3991\,
            in3 => \N__4005\,
            lcout => \o_LED_33_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_1_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4185\,
            in2 => \_gnd_net_\,
            in3 => \N__4209\,
            lcout => \r_count_5hzZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_2_c_RNO_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4168\,
            in1 => \N__4184\,
            in2 => \N__4150\,
            in3 => \N__4362\,
            lcout => \o_LED_23_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_3_c_RNO_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4303\,
            in1 => \N__4288\,
            in2 => \N__4348\,
            in3 => \N__4272\,
            lcout => \o_LED_23_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4208\,
            in2 => \_gnd_net_\,
            in3 => \N__3567\,
            lcout => \r_count_5hzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_7_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4312\,
            in1 => \_gnd_net_\,
            in2 => \N__3571\,
            in3 => \N__4330\,
            lcout => \r_count_5hzZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_12_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4572\,
            in1 => \N__4558\,
            in2 => \_gnd_net_\,
            in3 => \N__3558\,
            lcout => \r_count_5hzZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_15_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4489\,
            in1 => \_gnd_net_\,
            in2 => \N__3570\,
            in3 => \N__4503\,
            lcout => \r_count_5hzZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_14_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4533\,
            in1 => \N__4513\,
            in2 => \_gnd_net_\,
            in3 => \N__3559\,
            lcout => \r_count_5hzZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_1_c_RNO_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4480\,
            in1 => \N__4502\,
            in2 => \N__4210\,
            in3 => \N__4448\,
            lcout => \o_LED_23_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_4_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4387\,
            in1 => \N__4372\,
            in2 => \_gnd_net_\,
            in3 => \N__3563\,
            lcout => \r_count_5hzZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6501\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_0_c_RNO_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4329\,
            in1 => \N__4386\,
            in2 => \N__4534\,
            in3 => \N__4571\,
            lcout => \o_LED_23_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_7_c_RNO_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4734\,
            in1 => \N__4752\,
            in2 => \N__4789\,
            in3 => \N__4767\,
            lcout => \o_LED_23_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_16_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4459\,
            in2 => \N__3568\,
            in3 => \N__4479\,
            lcout => \r_count_5hzZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_5_c_RNO_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4704\,
            in1 => \N__4653\,
            in2 => \N__4672\,
            in3 => \N__4690\,
            lcout => \o_LED_23_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LEDZ0Z_2_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3569\,
            in3 => \N__3369\,
            lcout => \o_LED_2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_6_c_RNO_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4635\,
            in1 => \N__4620\,
            in2 => \N__4606\,
            in3 => \N__4587\,
            lcout => \o_LED_23_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_23_4_c_RNO_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4549\,
            in1 => \N__4258\,
            in2 => \N__4423\,
            in3 => \N__4401\,
            lcout => \o_LED_23_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_17_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4432\,
            in1 => \N__4450\,
            in2 => \_gnd_net_\,
            in3 => \N__3554\,
            lcout => \r_count_5hzZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_1_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3523\,
            in2 => \N__3505\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un2_r_count_2hz_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3483\,
            in2 => \_gnd_net_\,
            in3 => \N__3469\,
            lcout => \r_count_2hzZ0Z_2\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_1,
            carryout => un2_r_count_2hz_1_cry_2,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3466\,
            in2 => \_gnd_net_\,
            in3 => \N__3454\,
            lcout => \r_count_2hzZ0Z_3\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_2,
            carryout => un2_r_count_2hz_1_cry_3,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_3_THRU_LUT4_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3449\,
            in2 => \_gnd_net_\,
            in3 => \N__3430\,
            lcout => \un2_r_count_2hz_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_3,
            carryout => un2_r_count_2hz_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_5_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3426\,
            in2 => \_gnd_net_\,
            in3 => \N__3415\,
            lcout => \r_count_2hzZ0Z_5\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_4,
            carryout => un2_r_count_2hz_1_cry_5,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_6_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3765\,
            in2 => \_gnd_net_\,
            in3 => \N__3754\,
            lcout => \r_count_2hzZ0Z_6\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_5,
            carryout => un2_r_count_2hz_1_cry_6,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_7_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3747\,
            in2 => \_gnd_net_\,
            in3 => \N__3736\,
            lcout => \r_count_2hzZ0Z_7\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_6,
            carryout => un2_r_count_2hz_1_cry_7,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_8_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3733\,
            in2 => \_gnd_net_\,
            in3 => \N__3721\,
            lcout => \r_count_2hzZ0Z_8\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_7,
            carryout => un2_r_count_2hz_1_cry_8,
            clk => \N__6492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_8_THRU_LUT4_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3713\,
            in2 => \_gnd_net_\,
            in3 => \N__3694\,
            lcout => \un2_r_count_2hz_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => un2_r_count_2hz_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_9_THRU_LUT4_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3683\,
            in2 => \_gnd_net_\,
            in3 => \N__3661\,
            lcout => \un2_r_count_2hz_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_9,
            carryout => un2_r_count_2hz_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_10_THRU_LUT4_0_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3658\,
            in2 => \_gnd_net_\,
            in3 => \N__3637\,
            lcout => \un2_r_count_2hz_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_10,
            carryout => un2_r_count_2hz_1_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_11_THRU_LUT4_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3632\,
            in2 => \_gnd_net_\,
            in3 => \N__3607\,
            lcout => \un2_r_count_2hz_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_11,
            carryout => un2_r_count_2hz_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_13_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3603\,
            in2 => \_gnd_net_\,
            in3 => \N__3592\,
            lcout => \r_count_2hzZ0Z_13\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_12,
            carryout => un2_r_count_2hz_1_cry_13,
            clk => \N__6489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_13_THRU_LUT4_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3969\,
            in2 => \_gnd_net_\,
            in3 => \N__3946\,
            lcout => \un2_r_count_2hz_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_13,
            carryout => un2_r_count_2hz_1_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_15_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3942\,
            in2 => \_gnd_net_\,
            in3 => \N__3928\,
            lcout => \r_count_2hzZ0Z_15\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_14,
            carryout => un2_r_count_2hz_1_cry_15,
            clk => \N__6489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_15_THRU_LUT4_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3924\,
            in2 => \_gnd_net_\,
            in3 => \N__3898\,
            lcout => \un2_r_count_2hz_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_15,
            carryout => un2_r_count_2hz_1_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_16_THRU_LUT4_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3895\,
            in2 => \_gnd_net_\,
            in3 => \N__3868\,
            lcout => \un2_r_count_2hz_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => un2_r_count_2hz_1_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_17_THRU_LUT4_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3864\,
            in2 => \_gnd_net_\,
            in3 => \N__3841\,
            lcout => \un2_r_count_2hz_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_17,
            carryout => un2_r_count_2hz_1_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_18_THRU_LUT4_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3837\,
            in2 => \_gnd_net_\,
            in3 => \N__3811\,
            lcout => \un2_r_count_2hz_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_18,
            carryout => un2_r_count_2hz_1_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_19_THRU_LUT4_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3807\,
            in2 => \_gnd_net_\,
            in3 => \N__3784\,
            lcout => \un2_r_count_2hz_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_19,
            carryout => un2_r_count_2hz_1_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_21_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3781\,
            in2 => \_gnd_net_\,
            in3 => \N__3769\,
            lcout => \r_count_2hzZ0Z_21\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_20,
            carryout => un2_r_count_2hz_1_cry_21,
            clk => \N__6486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_2hz_1_cry_21_THRU_LUT4_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4130\,
            in2 => \_gnd_net_\,
            in3 => \N__4105\,
            lcout => \un2_r_count_2hz_1_cry_21_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_21,
            carryout => un2_r_count_2hz_1_cry_22,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_23_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4102\,
            in2 => \_gnd_net_\,
            in3 => \N__4090\,
            lcout => \r_count_2hzZ0Z_23\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_22,
            carryout => un2_r_count_2hz_1_cry_23,
            clk => \N__6486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_24_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4086\,
            in2 => \_gnd_net_\,
            in3 => \N__4072\,
            lcout => \r_count_2hzZ0Z_24\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_23,
            carryout => un2_r_count_2hz_1_cry_24,
            clk => \N__6486\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_25_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4069\,
            in2 => \_gnd_net_\,
            in3 => \N__4057\,
            lcout => \r_count_2hzZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => un2_r_count_2hz_1_cry_25,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_26_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4053\,
            in2 => \_gnd_net_\,
            in3 => \N__4039\,
            lcout => \r_count_2hzZ0Z_26\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_25,
            carryout => un2_r_count_2hz_1_cry_26,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_27_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4036\,
            in2 => \_gnd_net_\,
            in3 => \N__4024\,
            lcout => \r_count_2hzZ0Z_27\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_26,
            carryout => un2_r_count_2hz_1_cry_27,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_28_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4021\,
            in2 => \_gnd_net_\,
            in3 => \N__4009\,
            lcout => \r_count_2hzZ0Z_28\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_27,
            carryout => un2_r_count_2hz_1_cry_28,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_29_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4006\,
            in2 => \_gnd_net_\,
            in3 => \N__3994\,
            lcout => \r_count_2hzZ0Z_29\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_28,
            carryout => un2_r_count_2hz_1_cry_29,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_30_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3990\,
            in2 => \_gnd_net_\,
            in3 => \N__3976\,
            lcout => \r_count_2hzZ0Z_30\,
            ltout => OPEN,
            carryin => un2_r_count_2hz_1_cry_29,
            carryout => un2_r_count_2hz_1_cry_30,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_2hz_31_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4240\,
            in2 => \_gnd_net_\,
            in3 => \N__4243\,
            lcout => \r_count_2hzZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_5_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5001\,
            in1 => \N__4984\,
            in2 => \_gnd_net_\,
            in3 => \N__4868\,
            lcout => \r_count_1hzZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_3_c_RNO_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5092\,
            in1 => \N__5116\,
            in2 => \N__5065\,
            in3 => \N__5041\,
            lcout => \o_LED_43_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LEDZ0Z_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4876\,
            in3 => \N__4221\,
            lcout => \o_LED_4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_0_c_RNO_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5305\,
            in1 => \N__5000\,
            in2 => \N__5269\,
            in3 => \N__5225\,
            lcout => \o_LED_43_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5120\,
            in2 => \_gnd_net_\,
            in3 => \N__4872\,
            lcout => \r_count_1hzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_1_c_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4204\,
            in2 => \N__4186\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => un2_r_count_5hz_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_2_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4164\,
            in2 => \_gnd_net_\,
            in3 => \N__4153\,
            lcout => \r_count_5hzZ0Z_2\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_1,
            carryout => un2_r_count_5hz_1_cry_2,
            clk => \N__6509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_3_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4146\,
            in2 => \_gnd_net_\,
            in3 => \N__4135\,
            lcout => \r_count_5hzZ0Z_3\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_2,
            carryout => un2_r_count_5hz_1_cry_3,
            clk => \N__6509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_3_THRU_LUT4_0_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4385\,
            in2 => \_gnd_net_\,
            in3 => \N__4366\,
            lcout => \un2_r_count_5hz_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_3,
            carryout => un2_r_count_5hz_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_5_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4363\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \r_count_5hzZ0Z_5\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_4,
            carryout => un2_r_count_5hz_1_cry_5,
            clk => \N__6509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_6_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4344\,
            in2 => \_gnd_net_\,
            in3 => \N__4333\,
            lcout => \r_count_5hzZ0Z_6\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_5,
            carryout => un2_r_count_5hz_1_cry_6,
            clk => \N__6509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_6_THRU_LUT4_0_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4328\,
            in2 => \_gnd_net_\,
            in3 => \N__4306\,
            lcout => \un2_r_count_5hz_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_6,
            carryout => un2_r_count_5hz_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_8_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4302\,
            in2 => \_gnd_net_\,
            in3 => \N__4291\,
            lcout => \r_count_5hzZ0Z_8\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_7,
            carryout => un2_r_count_5hz_1_cry_8,
            clk => \N__6509\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_9_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4287\,
            in2 => \_gnd_net_\,
            in3 => \N__4276\,
            lcout => \r_count_5hzZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => un2_r_count_5hz_1_cry_9,
            clk => \N__6506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_10_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4273\,
            in2 => \_gnd_net_\,
            in3 => \N__4261\,
            lcout => \r_count_5hzZ0Z_10\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_9,
            carryout => un2_r_count_5hz_1_cry_10,
            clk => \N__6506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_11_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4257\,
            in2 => \_gnd_net_\,
            in3 => \N__4246\,
            lcout => \r_count_5hzZ0Z_11\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_10,
            carryout => un2_r_count_5hz_1_cry_11,
            clk => \N__6506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_11_THRU_LUT4_0_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4573\,
            in2 => \_gnd_net_\,
            in3 => \N__4552\,
            lcout => \un2_r_count_5hz_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_11,
            carryout => un2_r_count_5hz_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_13_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \N__4537\,
            lcout => \r_count_5hzZ0Z_13\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_12,
            carryout => un2_r_count_5hz_1_cry_13,
            clk => \N__6506\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_13_THRU_LUT4_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4532\,
            in2 => \_gnd_net_\,
            in3 => \N__4507\,
            lcout => \un2_r_count_5hz_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_13,
            carryout => un2_r_count_5hz_1_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_14_THRU_LUT4_0_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4504\,
            in2 => \_gnd_net_\,
            in3 => \N__4483\,
            lcout => \un2_r_count_5hz_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_14,
            carryout => un2_r_count_5hz_1_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_15_THRU_LUT4_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4478\,
            in2 => \_gnd_net_\,
            in3 => \N__4453\,
            lcout => \un2_r_count_5hz_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_15,
            carryout => un2_r_count_5hz_1_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_5hz_1_cry_16_THRU_LUT4_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4449\,
            in2 => \_gnd_net_\,
            in3 => \N__4426\,
            lcout => \un2_r_count_5hz_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => un2_r_count_5hz_1_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_18_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4422\,
            in2 => \_gnd_net_\,
            in3 => \N__4405\,
            lcout => \r_count_5hzZ0Z_18\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_17,
            carryout => un2_r_count_5hz_1_cry_18,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_19_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4402\,
            in2 => \_gnd_net_\,
            in3 => \N__4390\,
            lcout => \r_count_5hzZ0Z_19\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_18,
            carryout => un2_r_count_5hz_1_cry_19,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_20_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4705\,
            in2 => \_gnd_net_\,
            in3 => \N__4693\,
            lcout => \r_count_5hzZ0Z_20\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_19,
            carryout => un2_r_count_5hz_1_cry_20,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_21_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__4675\,
            lcout => \r_count_5hzZ0Z_21\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_20,
            carryout => un2_r_count_5hz_1_cry_21,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_22_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4671\,
            in2 => \_gnd_net_\,
            in3 => \N__4657\,
            lcout => \r_count_5hzZ0Z_22\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_21,
            carryout => un2_r_count_5hz_1_cry_22,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_23_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4654\,
            in2 => \_gnd_net_\,
            in3 => \N__4639\,
            lcout => \r_count_5hzZ0Z_23\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_22,
            carryout => un2_r_count_5hz_1_cry_23,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_24_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4636\,
            in2 => \_gnd_net_\,
            in3 => \N__4624\,
            lcout => \r_count_5hzZ0Z_24\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_23,
            carryout => un2_r_count_5hz_1_cry_24,
            clk => \N__6502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_25_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4621\,
            in2 => \_gnd_net_\,
            in3 => \N__4609\,
            lcout => \r_count_5hzZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => un2_r_count_5hz_1_cry_25,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_26_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4605\,
            in2 => \_gnd_net_\,
            in3 => \N__4591\,
            lcout => \r_count_5hzZ0Z_26\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_25,
            carryout => un2_r_count_5hz_1_cry_26,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_27_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4588\,
            in2 => \_gnd_net_\,
            in3 => \N__4576\,
            lcout => \r_count_5hzZ0Z_27\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_26,
            carryout => un2_r_count_5hz_1_cry_27,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_28_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4785\,
            in2 => \_gnd_net_\,
            in3 => \N__4771\,
            lcout => \r_count_5hzZ0Z_28\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_27,
            carryout => un2_r_count_5hz_1_cry_28,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_29_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4768\,
            in2 => \_gnd_net_\,
            in3 => \N__4756\,
            lcout => \r_count_5hzZ0Z_29\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_28,
            carryout => un2_r_count_5hz_1_cry_29,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_30_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4753\,
            in2 => \_gnd_net_\,
            in3 => \N__4741\,
            lcout => \r_count_5hzZ0Z_30\,
            ltout => OPEN,
            carryin => un2_r_count_5hz_1_cry_29,
            carryout => un2_r_count_5hz_1_cry_30,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_5hz_31_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4735\,
            in2 => \_gnd_net_\,
            in3 => \N__4738\,
            lcout => \r_count_5hzZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_0_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4723\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \o_LED_43_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_1_c_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4807\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_0\,
            carryout => \o_LED_43_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_2_c_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4798\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_1\,
            carryout => \o_LED_43_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_3_c_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4714\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_2\,
            carryout => \o_LED_43_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_4_c_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5143\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_3\,
            carryout => \o_LED_43_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_5_c_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6364\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_4\,
            carryout => \o_LED_43_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_6_c_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_5\,
            carryout => \o_LED_43_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_7_c_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5740\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_43_6\,
            carryout => \o_LED_43\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_THRU_LUT4_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4813\,
            lcout => \o_LED_43_THRU_CO\,
            ltout => \o_LED_43_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_15_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5161\,
            in2 => \N__4810\,
            in3 => \N__5572\,
            lcout => \r_count_1hzZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_1_c_RNO_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5160\,
            in1 => \N__5192\,
            in2 => \N__5556\,
            in3 => \N__5510\,
            lcout => \o_LED_43_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_10_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5284\,
            in1 => \N__5303\,
            in2 => \_gnd_net_\,
            in3 => \N__4852\,
            lcout => \r_count_1hzZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_2_c_RNO_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5373\,
            in1 => \N__5441\,
            in2 => \N__5412\,
            in3 => \N__5477\,
            lcout => \o_LED_43_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_12_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5209\,
            in1 => \N__5229\,
            in2 => \_gnd_net_\,
            in3 => \N__4854\,
            lcout => \r_count_1hzZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_13_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5176\,
            in1 => \_gnd_net_\,
            in2 => \N__4873\,
            in3 => \N__5193\,
            lcout => \r_count_1hzZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_11_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5245\,
            in1 => \N__5267\,
            in2 => \_gnd_net_\,
            in3 => \N__4853\,
            lcout => \r_count_1hzZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_23_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__5372\,
            in2 => \_gnd_net_\,
            in3 => \N__4867\,
            lcout => \r_count_1hzZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_21_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5389\,
            in2 => \N__4875\,
            in3 => \N__5411\,
            lcout => \r_count_1hzZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_18_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5497\,
            in1 => \N__5518\,
            in2 => \_gnd_net_\,
            in3 => \N__4859\,
            lcout => \r_count_1hzZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_20_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5425\,
            in1 => \N__5445\,
            in2 => \_gnd_net_\,
            in3 => \N__4863\,
            lcout => \r_count_1hzZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_19_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5461\,
            in2 => \N__4874\,
            in3 => \N__5481\,
            lcout => \r_count_1hzZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_17_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5533\,
            in1 => \N__5555\,
            in2 => \_gnd_net_\,
            in3 => \N__4858\,
            lcout => \r_count_1hzZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_0_c_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5677\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_1_0_\,
            carryout => \o_LED_13_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_1_c_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_0\,
            carryout => \o_LED_13_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_2_c_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5659\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_1\,
            carryout => \o_LED_13_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_3_c_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5668\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_2\,
            carryout => \o_LED_13_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_4_c_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4936\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_3\,
            carryout => \o_LED_13_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_5_c_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4924\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_4\,
            carryout => \o_LED_13_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_6_c_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_5\,
            carryout => \o_LED_13_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_7_c_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4903\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \o_LED_13_6\,
            carryout => \o_LED_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_THRU_LUT4_0_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4891\,
            lcout => \o_LED_13_THRU_CO\,
            ltout => \o_LED_13_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_4_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5911\,
            in2 => \N__4888\,
            in3 => \N__5929\,
            lcout => \r_count_10hzZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6512\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_1_c_RNO_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6035\,
            in1 => \N__6005\,
            in2 => \N__6112\,
            in3 => \N__6263\,
            lcout => \o_LED_13_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_20_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6247\,
            in2 => \N__5724\,
            in3 => \N__6267\,
            lcout => \r_count_10hzZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_12_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6091\,
            in2 => \N__5721\,
            in3 => \N__6111\,
            lcout => \r_count_10hzZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LEDZ0Z_1_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4947\,
            in2 => \_gnd_net_\,
            in3 => \N__5715\,
            lcout => \o_LED_1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_17_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5989\,
            in2 => \N__5723\,
            in3 => \N__6009\,
            lcout => \r_count_10hzZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_9_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5800\,
            in1 => \N__5818\,
            in2 => \_gnd_net_\,
            in3 => \N__5714\,
            lcout => \r_count_10hzZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_16_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6019\,
            in2 => \N__5722\,
            in3 => \N__6037\,
            lcout => \r_count_10hzZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_4_c_RNO_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__6066\,
            in2 => \N__5977\,
            in3 => \N__6081\,
            lcout => \o_LED_13_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_5_c_RNO_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6195\,
            in1 => \N__6235\,
            in2 => \N__6217\,
            in3 => \N__6285\,
            lcout => \o_LED_13_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_6_c_RNO_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6180\,
            in1 => \N__6591\,
            in2 => \N__6166\,
            in3 => \N__6147\,
            lcout => \o_LED_13_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_7_c_RNO_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6543\,
            in1 => \N__6525\,
            in2 => \N__6577\,
            in3 => \N__6558\,
            lcout => \o_LED_13_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5087\,
            in2 => \_gnd_net_\,
            in3 => \N__5128\,
            lcout => \r_count_1hzZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6493\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_4_c_RNO_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4969\,
            in1 => \N__5020\,
            in2 => \N__5341\,
            in3 => \N__5322\,
            lcout => \o_LED_43_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_1_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5127\,
            in2 => \N__5088\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => un2_r_count_1hz_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5055\,
            in2 => \_gnd_net_\,
            in3 => \N__5044\,
            lcout => \r_count_1hzZ0Z_2\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_1,
            carryout => un2_r_count_1hz_1_cry_2,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5037\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \r_count_1hzZ0Z_3\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_2,
            carryout => un2_r_count_1hz_1_cry_3,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5019\,
            in2 => \_gnd_net_\,
            in3 => \N__5008\,
            lcout => \r_count_1hzZ0Z_4\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_3,
            carryout => un2_r_count_1hz_1_cry_4,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_4_THRU_LUT4_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5005\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => \un2_r_count_1hz_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_4,
            carryout => un2_r_count_1hz_1_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4968\,
            in2 => \_gnd_net_\,
            in3 => \N__4957\,
            lcout => \r_count_1hzZ0Z_6\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_5,
            carryout => un2_r_count_1hz_1_cry_6,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5337\,
            in2 => \_gnd_net_\,
            in3 => \N__5326\,
            lcout => \r_count_1hzZ0Z_7\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_6,
            carryout => un2_r_count_1hz_1_cry_7,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5323\,
            in2 => \_gnd_net_\,
            in3 => \N__5311\,
            lcout => \r_count_1hzZ0Z_8\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_7,
            carryout => un2_r_count_1hz_1_cry_8,
            clk => \N__6496\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_9_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6390\,
            in2 => \_gnd_net_\,
            in3 => \N__5308\,
            lcout => \r_count_1hzZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => un2_r_count_1hz_1_cry_9,
            clk => \N__6500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_9_THRU_LUT4_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5304\,
            in2 => \_gnd_net_\,
            in3 => \N__5272\,
            lcout => \un2_r_count_1hz_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_9,
            carryout => un2_r_count_1hz_1_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_10_THRU_LUT4_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5268\,
            in2 => \_gnd_net_\,
            in3 => \N__5233\,
            lcout => \un2_r_count_1hz_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_10,
            carryout => un2_r_count_1hz_1_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_11_THRU_LUT4_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5230\,
            in2 => \_gnd_net_\,
            in3 => \N__5197\,
            lcout => \un2_r_count_1hz_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_11,
            carryout => un2_r_count_1hz_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_12_THRU_LUT4_0_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5194\,
            in2 => \_gnd_net_\,
            in3 => \N__5167\,
            lcout => \un2_r_count_1hz_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_12,
            carryout => un2_r_count_1hz_1_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_14_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6415\,
            in2 => \_gnd_net_\,
            in3 => \N__5164\,
            lcout => \r_count_1hzZ0Z_14\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_13,
            carryout => un2_r_count_1hz_1_cry_14,
            clk => \N__6500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_14_THRU_LUT4_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5159\,
            in2 => \_gnd_net_\,
            in3 => \N__5563\,
            lcout => \un2_r_count_1hz_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_14,
            carryout => un2_r_count_1hz_1_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_16_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6376\,
            in2 => \_gnd_net_\,
            in3 => \N__5560\,
            lcout => \r_count_1hzZ0Z_16\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_15,
            carryout => un2_r_count_1hz_1_cry_16,
            clk => \N__6500\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_16_THRU_LUT4_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5557\,
            in2 => \_gnd_net_\,
            in3 => \N__5521\,
            lcout => \un2_r_count_1hz_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => un2_r_count_1hz_1_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_17_THRU_LUT4_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5517\,
            in2 => \_gnd_net_\,
            in3 => \N__5485\,
            lcout => \un2_r_count_1hz_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_17,
            carryout => un2_r_count_1hz_1_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_18_THRU_LUT4_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5482\,
            in2 => \_gnd_net_\,
            in3 => \N__5449\,
            lcout => \un2_r_count_1hz_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_18,
            carryout => un2_r_count_1hz_1_cry_19,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_19_THRU_LUT4_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5446\,
            in2 => \_gnd_net_\,
            in3 => \N__5416\,
            lcout => \un2_r_count_1hz_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_19,
            carryout => un2_r_count_1hz_1_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_20_THRU_LUT4_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5413\,
            in2 => \_gnd_net_\,
            in3 => \N__5380\,
            lcout => \un2_r_count_1hz_1_cry_20_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_20,
            carryout => un2_r_count_1hz_1_cry_21,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_22_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6403\,
            in2 => \_gnd_net_\,
            in3 => \N__5377\,
            lcout => \r_count_1hzZ0Z_22\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_21,
            carryout => un2_r_count_1hz_1_cry_22,
            clk => \N__6503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_1hz_1_cry_22_THRU_LUT4_0_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5374\,
            in2 => \_gnd_net_\,
            in3 => \N__5608\,
            lcout => \un2_r_count_1hz_1_cry_22_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_22,
            carryout => un2_r_count_1hz_1_cry_23,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_24_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6327\,
            in2 => \_gnd_net_\,
            in3 => \N__5605\,
            lcout => \r_count_1hzZ0Z_24\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_23,
            carryout => un2_r_count_1hz_1_cry_24,
            clk => \N__6503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_25_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6352\,
            in2 => \_gnd_net_\,
            in3 => \N__5602\,
            lcout => \r_count_1hzZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => un2_r_count_1hz_1_cry_25,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_26_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6340\,
            in2 => \_gnd_net_\,
            in3 => \N__5599\,
            lcout => \r_count_1hzZ0Z_26\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_25,
            carryout => un2_r_count_1hz_1_cry_26,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_27_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6313\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => \r_count_1hzZ0Z_27\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_26,
            carryout => un2_r_count_1hz_1_cry_27,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_28_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5764\,
            in3 => \N__5593\,
            lcout => \r_count_1hzZ0Z_28\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_27,
            carryout => un2_r_count_1hz_1_cry_28,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_29_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5581\,
            in2 => \_gnd_net_\,
            in3 => \N__5590\,
            lcout => \r_count_1hzZ0Z_29\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_28,
            carryout => un2_r_count_1hz_1_cry_29,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_30_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5749\,
            in2 => \_gnd_net_\,
            in3 => \N__5587\,
            lcout => \r_count_1hzZ0Z_30\,
            ltout => OPEN,
            carryin => un2_r_count_1hz_1_cry_29,
            carryout => un2_r_count_1hz_1_cry_30,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_1hz_31_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5773\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5584\,
            lcout => \r_count_1hzZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_7_c_RNO_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5580\,
            in1 => \N__5772\,
            in2 => \N__5763\,
            in3 => \N__5748\,
            lcout => \o_LED_43_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_6_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5887\,
            in1 => \N__5869\,
            in2 => \_gnd_net_\,
            in3 => \N__5716\,
            lcout => \r_count_10hzZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_7_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__5859\,
            in1 => \N__5842\,
            in2 => \N__5725\,
            in3 => \_gnd_net_\,
            lcout => \r_count_10hzZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_0_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5720\,
            lcout => \r_count_10hzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_0_c_RNO_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__5928\,
            in2 => \N__5860\,
            in3 => \N__5816\,
            lcout => \o_LED_13_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_1_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5629\,
            in1 => \_gnd_net_\,
            in2 => \N__5653\,
            in3 => \_gnd_net_\,
            lcout => \r_count_10hzZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6514\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_3_c_RNO_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5833\,
            in1 => \N__5902\,
            in2 => \N__5791\,
            in3 => \N__6130\,
            lcout => \o_LED_13_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_13_2_c_RNO_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5628\,
            in1 => \N__5959\,
            in2 => \N__5652\,
            in3 => \N__5943\,
            lcout => \o_LED_13_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_1_c_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5644\,
            in2 => \N__5627\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => un2_r_count_10hz_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5958\,
            in2 => \_gnd_net_\,
            in3 => \N__5947\,
            lcout => \r_count_10hzZ0Z_2\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_1,
            carryout => un2_r_count_10hz_1_cry_2,
            clk => \N__6513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_3_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5944\,
            in2 => \_gnd_net_\,
            in3 => \N__5932\,
            lcout => \r_count_10hzZ0Z_3\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_2,
            carryout => un2_r_count_10hz_1_cry_3,
            clk => \N__6513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_3_THRU_LUT4_0_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5927\,
            in2 => \_gnd_net_\,
            in3 => \N__5905\,
            lcout => \un2_r_count_10hz_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_3,
            carryout => un2_r_count_10hz_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_5_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5901\,
            in2 => \_gnd_net_\,
            in3 => \N__5890\,
            lcout => \r_count_10hzZ0Z_5\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_4,
            carryout => un2_r_count_10hz_1_cry_5,
            clk => \N__6513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_5_THRU_LUT4_0_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5885\,
            in2 => \_gnd_net_\,
            in3 => \N__5863\,
            lcout => \un2_r_count_10hz_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_5,
            carryout => un2_r_count_10hz_1_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_6_THRU_LUT4_0_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5855\,
            in2 => \_gnd_net_\,
            in3 => \N__5836\,
            lcout => \un2_r_count_10hz_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_6,
            carryout => un2_r_count_10hz_1_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_8_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5832\,
            in2 => \_gnd_net_\,
            in3 => \N__5821\,
            lcout => \r_count_10hzZ0Z_8\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_7,
            carryout => un2_r_count_10hz_1_cry_8,
            clk => \N__6513\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_8_THRU_LUT4_0_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5817\,
            in2 => \_gnd_net_\,
            in3 => \N__5794\,
            lcout => \un2_r_count_10hz_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => un2_r_count_10hz_1_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_10_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5787\,
            in2 => \_gnd_net_\,
            in3 => \N__6133\,
            lcout => \r_count_10hzZ0Z_10\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_9,
            carryout => un2_r_count_10hz_1_cry_10,
            clk => \N__6511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_11_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6129\,
            in2 => \_gnd_net_\,
            in3 => \N__6115\,
            lcout => \r_count_10hzZ0Z_11\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_10,
            carryout => un2_r_count_10hz_1_cry_11,
            clk => \N__6511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_11_THRU_LUT4_0_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6110\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => \un2_r_count_10hz_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_11,
            carryout => un2_r_count_10hz_1_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_13_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6082\,
            in2 => \_gnd_net_\,
            in3 => \N__6070\,
            lcout => \r_count_10hzZ0Z_13\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_12,
            carryout => un2_r_count_10hz_1_cry_13,
            clk => \N__6511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_14_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6067\,
            in2 => \_gnd_net_\,
            in3 => \N__6055\,
            lcout => \r_count_10hzZ0Z_14\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_13,
            carryout => un2_r_count_10hz_1_cry_14,
            clk => \N__6511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_15_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6052\,
            in2 => \_gnd_net_\,
            in3 => \N__6040\,
            lcout => \r_count_10hzZ0Z_15\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_14,
            carryout => un2_r_count_10hz_1_cry_15,
            clk => \N__6511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_15_THRU_LUT4_0_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6036\,
            in2 => \_gnd_net_\,
            in3 => \N__6013\,
            lcout => \un2_r_count_10hz_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_15,
            carryout => un2_r_count_10hz_1_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_16_THRU_LUT4_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6010\,
            in2 => \_gnd_net_\,
            in3 => \N__5980\,
            lcout => \un2_r_count_10hz_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => un2_r_count_10hz_1_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_18_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5976\,
            in2 => \_gnd_net_\,
            in3 => \N__5962\,
            lcout => \r_count_10hzZ0Z_18\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_17,
            carryout => un2_r_count_10hz_1_cry_18,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_19_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6286\,
            in2 => \_gnd_net_\,
            in3 => \N__6271\,
            lcout => \r_count_10hzZ0Z_19\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_18,
            carryout => un2_r_count_10hz_1_cry_19,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un2_r_count_10hz_1_cry_19_THRU_LUT4_0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6268\,
            in2 => \_gnd_net_\,
            in3 => \N__6238\,
            lcout => \un2_r_count_10hz_1_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_19,
            carryout => un2_r_count_10hz_1_cry_20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_21_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6234\,
            in2 => \_gnd_net_\,
            in3 => \N__6220\,
            lcout => \r_count_10hzZ0Z_21\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_20,
            carryout => un2_r_count_10hz_1_cry_21,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_22_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6213\,
            in2 => \_gnd_net_\,
            in3 => \N__6199\,
            lcout => \r_count_10hzZ0Z_22\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_21,
            carryout => un2_r_count_10hz_1_cry_22,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_23_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6196\,
            in2 => \_gnd_net_\,
            in3 => \N__6184\,
            lcout => \r_count_10hzZ0Z_23\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_22,
            carryout => un2_r_count_10hz_1_cry_23,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_24_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6181\,
            in2 => \_gnd_net_\,
            in3 => \N__6169\,
            lcout => \r_count_10hzZ0Z_24\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_23,
            carryout => un2_r_count_10hz_1_cry_24,
            clk => \N__6508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_25_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6165\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \r_count_10hzZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => un2_r_count_10hz_1_cry_25,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_26_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6148\,
            in2 => \_gnd_net_\,
            in3 => \N__6136\,
            lcout => \r_count_10hzZ0Z_26\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_25,
            carryout => un2_r_count_10hz_1_cry_26,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_27_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6592\,
            in2 => \_gnd_net_\,
            in3 => \N__6580\,
            lcout => \r_count_10hzZ0Z_27\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_26,
            carryout => un2_r_count_10hz_1_cry_27,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_28_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6576\,
            in2 => \_gnd_net_\,
            in3 => \N__6562\,
            lcout => \r_count_10hzZ0Z_28\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_27,
            carryout => un2_r_count_10hz_1_cry_28,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_29_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6559\,
            in2 => \_gnd_net_\,
            in3 => \N__6547\,
            lcout => \r_count_10hzZ0Z_29\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_28,
            carryout => un2_r_count_10hz_1_cry_29,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_30_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6544\,
            in2 => \_gnd_net_\,
            in3 => \N__6532\,
            lcout => \r_count_10hzZ0Z_30\,
            ltout => OPEN,
            carryin => un2_r_count_10hz_1_cry_29,
            carryout => un2_r_count_10hz_1_cry_30,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \r_count_10hz_31_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6526\,
            in2 => \_gnd_net_\,
            in3 => \N__6529\,
            lcout => \r_count_10hzZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_5_c_RNO_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6414\,
            in1 => \N__6402\,
            in2 => \N__6391\,
            in3 => \N__6375\,
            lcout => \o_LED_43_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_LED_43_6_c_RNO_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6351\,
            in1 => \N__6339\,
            in2 => \N__6328\,
            in3 => \N__6312\,
            lcout => \o_LED_43_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
