// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Oct 8 2022 16:56:32

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "LED_blink" view "INTERFACE"

module LED_blink (
    o_LED_3,
    o_LED_1,
    i_Clk,
    o_LED_4,
    o_LED_2);

    output o_LED_3;
    output o_LED_1;
    input i_Clk;
    output o_LED_4;
    output o_LED_2;

    wire N__6649;
    wire N__6648;
    wire N__6647;
    wire N__6638;
    wire N__6637;
    wire N__6636;
    wire N__6629;
    wire N__6628;
    wire N__6627;
    wire N__6620;
    wire N__6619;
    wire N__6618;
    wire N__6611;
    wire N__6610;
    wire N__6609;
    wire N__6592;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6580;
    wire N__6577;
    wire N__6576;
    wire N__6573;
    wire N__6570;
    wire N__6567;
    wire N__6562;
    wire N__6559;
    wire N__6558;
    wire N__6555;
    wire N__6552;
    wire N__6547;
    wire N__6544;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6514;
    wire N__6513;
    wire N__6512;
    wire N__6511;
    wire N__6510;
    wire N__6509;
    wire N__6508;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6504;
    wire N__6503;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6490;
    wire N__6489;
    wire N__6488;
    wire N__6487;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6403;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6376;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6340;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6328;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6267;
    wire N__6264;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6184;
    wire N__6181;
    wire N__6180;
    wire N__6177;
    wire N__6174;
    wire N__6169;
    wire N__6166;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6151;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6115;
    wire N__6112;
    wire N__6111;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6070;
    wire N__6067;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6055;
    wire N__6052;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6009;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5947;
    wire N__5944;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5932;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5890;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5859;
    wire N__5856;
    wire N__5855;
    wire N__5850;
    wire N__5847;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5821;
    wire N__5818;
    wire N__5817;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5773;
    wire N__5772;
    wire N__5767;
    wire N__5764;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5752;
    wire N__5749;
    wire N__5748;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5724;
    wire N__5723;
    wire N__5722;
    wire N__5721;
    wire N__5720;
    wire N__5717;
    wire N__5716;
    wire N__5715;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5695;
    wire N__5682;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5652;
    wire N__5649;
    wire N__5648;
    wire N__5645;
    wire N__5644;
    wire N__5637;
    wire N__5634;
    wire N__5629;
    wire N__5628;
    wire N__5627;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5613;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5580;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5510;
    wire N__5505;
    wire N__5502;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5481;
    wire N__5478;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5445;
    wire N__5442;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5412;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5373;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5326;
    wire N__5323;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5304;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5289;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5268;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5229;
    wire N__5226;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5216;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5184;
    wire N__5181;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5160;
    wire N__5159;
    wire N__5154;
    wire N__5151;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5120;
    wire N__5117;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5055;
    wire N__5052;
    wire N__5049;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5023;
    wire N__5020;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__5001;
    wire N__5000;
    wire N__4997;
    wire N__4992;
    wire N__4989;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4957;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4876;
    wire N__4875;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4869;
    wire N__4868;
    wire N__4867;
    wire N__4864;
    wire N__4863;
    wire N__4860;
    wire N__4859;
    wire N__4858;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4844;
    wire N__4831;
    wire N__4822;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4771;
    wire N__4768;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4756;
    wire N__4753;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4734;
    wire N__4731;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4675;
    wire N__4672;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4624;
    wire N__4621;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4609;
    wire N__4606;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4591;
    wire N__4588;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4576;
    wire N__4573;
    wire N__4572;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4537;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4503;
    wire N__4502;
    wire N__4499;
    wire N__4494;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4479;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4449;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4422;
    wire N__4419;
    wire N__4416;
    wire N__4413;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4401;
    wire N__4398;
    wire N__4395;
    wire N__4390;
    wire N__4387;
    wire N__4386;
    wire N__4385;
    wire N__4380;
    wire N__4377;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4333;
    wire N__4330;
    wire N__4329;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4291;
    wire N__4288;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4276;
    wire N__4273;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4210;
    wire N__4209;
    wire N__4208;
    wire N__4205;
    wire N__4204;
    wire N__4201;
    wire N__4196;
    wire N__4193;
    wire N__4186;
    wire N__4185;
    wire N__4184;
    wire N__4181;
    wire N__4176;
    wire N__4173;
    wire N__4168;
    wire N__4165;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4135;
    wire N__4132;
    wire N__4131;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4090;
    wire N__4087;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4072;
    wire N__4069;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4057;
    wire N__4054;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4039;
    wire N__4036;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4024;
    wire N__4021;
    wire N__4020;
    wire N__4017;
    wire N__4014;
    wire N__4009;
    wire N__4006;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3994;
    wire N__3991;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3969;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3933;
    wire N__3928;
    wire N__3925;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3891;
    wire N__3890;
    wire N__3887;
    wire N__3882;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3864;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3837;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3807;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3769;
    wire N__3766;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3736;
    wire N__3733;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3714;
    wire N__3713;
    wire N__3708;
    wire N__3705;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3690;
    wire N__3687;
    wire N__3684;
    wire N__3683;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3657;
    wire N__3656;
    wire N__3653;
    wire N__3648;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3633;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3592;
    wire N__3589;
    wire N__3586;
    wire N__3583;
    wire N__3580;
    wire N__3577;
    wire N__3574;
    wire N__3571;
    wire N__3570;
    wire N__3569;
    wire N__3568;
    wire N__3567;
    wire N__3564;
    wire N__3563;
    wire N__3560;
    wire N__3559;
    wire N__3558;
    wire N__3555;
    wire N__3554;
    wire N__3551;
    wire N__3538;
    wire N__3531;
    wire N__3526;
    wire N__3525;
    wire N__3524;
    wire N__3523;
    wire N__3520;
    wire N__3515;
    wire N__3512;
    wire N__3505;
    wire N__3504;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3491;
    wire N__3484;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3469;
    wire N__3466;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3454;
    wire N__3451;
    wire N__3450;
    wire N__3449;
    wire N__3444;
    wire N__3441;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3358;
    wire N__3357;
    wire N__3356;
    wire N__3355;
    wire N__3354;
    wire N__3353;
    wire N__3352;
    wire N__3349;
    wire N__3348;
    wire N__3345;
    wire N__3342;
    wire N__3341;
    wire N__3338;
    wire N__3337;
    wire N__3336;
    wire N__3333;
    wire N__3332;
    wire N__3329;
    wire N__3328;
    wire N__3325;
    wire N__3314;
    wire N__3299;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire N__3223;
    wire N__3220;
    wire N__3217;
    wire N__3214;
    wire N__3211;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3198;
    wire N__3195;
    wire N__3192;
    wire N__3187;
    wire N__3184;
    wire N__3181;
    wire N__3178;
    wire N__3175;
    wire N__3172;
    wire VCCG0;
    wire GNDG0;
    wire bfn_6_7_0_;
    wire o_LED_33_0;
    wire o_LED_33_1;
    wire o_LED_33_2;
    wire o_LED_33_3;
    wire o_LED_33_4;
    wire o_LED_33_5;
    wire o_LED_33_6;
    wire o_LED_33;
    wire bfn_6_8_0_;
    wire o_LED_33_THRU_CO_cascade_;
    wire o_LED_3_c;
    wire o_LED_33_2_and;
    wire o_LED_33_1_and;
    wire bfn_7_3_0_;
    wire o_LED_23_0;
    wire o_LED_23_1;
    wire o_LED_23_2;
    wire o_LED_23_3;
    wire o_LED_23_4;
    wire o_LED_23_5;
    wire o_LED_23_6;
    wire o_LED_23;
    wire bfn_7_4_0_;
    wire o_LED_33_4_and;
    wire o_LED_33_3_and;
    wire o_LED_33_5_and;
    wire o_LED_33_0_and;
    wire o_LED_33_6_and;
    wire o_LED_33_THRU_CO;
    wire o_LED_33_7_and;
    wire o_LED_23_2_and;
    wire o_LED_23_3_and;
    wire o_LED_23_1_and;
    wire o_LED_23_0_and;
    wire o_LED_23_7_and;
    wire o_LED_23_5_and;
    wire o_LED_2_c;
    wire o_LED_23_6_and;
    wire o_LED_23_4_and;
    wire o_LED_23_THRU_CO;
    wire r_count_2hzZ0Z_0;
    wire r_count_2hzZ0Z_1;
    wire bfn_8_6_0_;
    wire r_count_2hzZ0Z_2;
    wire un2_r_count_2hz_1_cry_1;
    wire r_count_2hzZ0Z_3;
    wire un2_r_count_2hz_1_cry_2;
    wire r_count_2hzZ0Z_4;
    wire un2_r_count_2hz_1_cry_3_THRU_CO;
    wire un2_r_count_2hz_1_cry_3;
    wire r_count_2hzZ0Z_5;
    wire un2_r_count_2hz_1_cry_4;
    wire r_count_2hzZ0Z_6;
    wire un2_r_count_2hz_1_cry_5;
    wire r_count_2hzZ0Z_7;
    wire un2_r_count_2hz_1_cry_6;
    wire r_count_2hzZ0Z_8;
    wire un2_r_count_2hz_1_cry_7;
    wire un2_r_count_2hz_1_cry_8;
    wire r_count_2hzZ0Z_9;
    wire un2_r_count_2hz_1_cry_8_THRU_CO;
    wire bfn_8_7_0_;
    wire r_count_2hzZ0Z_10;
    wire un2_r_count_2hz_1_cry_9_THRU_CO;
    wire un2_r_count_2hz_1_cry_9;
    wire r_count_2hzZ0Z_11;
    wire un2_r_count_2hz_1_cry_10_THRU_CO;
    wire un2_r_count_2hz_1_cry_10;
    wire r_count_2hzZ0Z_12;
    wire un2_r_count_2hz_1_cry_11_THRU_CO;
    wire un2_r_count_2hz_1_cry_11;
    wire r_count_2hzZ0Z_13;
    wire un2_r_count_2hz_1_cry_12;
    wire r_count_2hzZ0Z_14;
    wire un2_r_count_2hz_1_cry_13_THRU_CO;
    wire un2_r_count_2hz_1_cry_13;
    wire r_count_2hzZ0Z_15;
    wire un2_r_count_2hz_1_cry_14;
    wire r_count_2hzZ0Z_16;
    wire un2_r_count_2hz_1_cry_15_THRU_CO;
    wire un2_r_count_2hz_1_cry_15;
    wire un2_r_count_2hz_1_cry_16;
    wire r_count_2hzZ0Z_17;
    wire un2_r_count_2hz_1_cry_16_THRU_CO;
    wire bfn_8_8_0_;
    wire r_count_2hzZ0Z_18;
    wire un2_r_count_2hz_1_cry_17_THRU_CO;
    wire un2_r_count_2hz_1_cry_17;
    wire r_count_2hzZ0Z_19;
    wire un2_r_count_2hz_1_cry_18_THRU_CO;
    wire un2_r_count_2hz_1_cry_18;
    wire r_count_2hzZ0Z_20;
    wire un2_r_count_2hz_1_cry_19_THRU_CO;
    wire un2_r_count_2hz_1_cry_19;
    wire r_count_2hzZ0Z_21;
    wire un2_r_count_2hz_1_cry_20;
    wire r_count_2hzZ0Z_22;
    wire un2_r_count_2hz_1_cry_21_THRU_CO;
    wire un2_r_count_2hz_1_cry_21;
    wire r_count_2hzZ0Z_23;
    wire un2_r_count_2hz_1_cry_22;
    wire r_count_2hzZ0Z_24;
    wire un2_r_count_2hz_1_cry_23;
    wire un2_r_count_2hz_1_cry_24;
    wire r_count_2hzZ0Z_25;
    wire bfn_8_9_0_;
    wire r_count_2hzZ0Z_26;
    wire un2_r_count_2hz_1_cry_25;
    wire r_count_2hzZ0Z_27;
    wire un2_r_count_2hz_1_cry_26;
    wire r_count_2hzZ0Z_28;
    wire un2_r_count_2hz_1_cry_27;
    wire r_count_2hzZ0Z_29;
    wire un2_r_count_2hz_1_cry_28;
    wire r_count_2hzZ0Z_30;
    wire un2_r_count_2hz_1_cry_29;
    wire un2_r_count_2hz_1_cry_30;
    wire r_count_2hzZ0Z_31;
    wire o_LED_4_c;
    wire r_count_5hzZ0Z_0;
    wire r_count_5hzZ0Z_1;
    wire bfn_9_2_0_;
    wire r_count_5hzZ0Z_2;
    wire un2_r_count_5hz_1_cry_1;
    wire r_count_5hzZ0Z_3;
    wire un2_r_count_5hz_1_cry_2;
    wire r_count_5hzZ0Z_4;
    wire un2_r_count_5hz_1_cry_3_THRU_CO;
    wire un2_r_count_5hz_1_cry_3;
    wire r_count_5hzZ0Z_5;
    wire un2_r_count_5hz_1_cry_4;
    wire r_count_5hzZ0Z_6;
    wire un2_r_count_5hz_1_cry_5;
    wire r_count_5hzZ0Z_7;
    wire un2_r_count_5hz_1_cry_6_THRU_CO;
    wire un2_r_count_5hz_1_cry_6;
    wire r_count_5hzZ0Z_8;
    wire un2_r_count_5hz_1_cry_7;
    wire un2_r_count_5hz_1_cry_8;
    wire r_count_5hzZ0Z_9;
    wire bfn_9_3_0_;
    wire r_count_5hzZ0Z_10;
    wire un2_r_count_5hz_1_cry_9;
    wire r_count_5hzZ0Z_11;
    wire un2_r_count_5hz_1_cry_10;
    wire r_count_5hzZ0Z_12;
    wire un2_r_count_5hz_1_cry_11_THRU_CO;
    wire un2_r_count_5hz_1_cry_11;
    wire r_count_5hzZ0Z_13;
    wire un2_r_count_5hz_1_cry_12;
    wire r_count_5hzZ0Z_14;
    wire un2_r_count_5hz_1_cry_13_THRU_CO;
    wire un2_r_count_5hz_1_cry_13;
    wire r_count_5hzZ0Z_15;
    wire un2_r_count_5hz_1_cry_14_THRU_CO;
    wire un2_r_count_5hz_1_cry_14;
    wire r_count_5hzZ0Z_16;
    wire un2_r_count_5hz_1_cry_15_THRU_CO;
    wire un2_r_count_5hz_1_cry_15;
    wire un2_r_count_5hz_1_cry_16;
    wire r_count_5hzZ0Z_17;
    wire un2_r_count_5hz_1_cry_16_THRU_CO;
    wire bfn_9_4_0_;
    wire r_count_5hzZ0Z_18;
    wire un2_r_count_5hz_1_cry_17;
    wire r_count_5hzZ0Z_19;
    wire un2_r_count_5hz_1_cry_18;
    wire r_count_5hzZ0Z_20;
    wire un2_r_count_5hz_1_cry_19;
    wire r_count_5hzZ0Z_21;
    wire un2_r_count_5hz_1_cry_20;
    wire r_count_5hzZ0Z_22;
    wire un2_r_count_5hz_1_cry_21;
    wire r_count_5hzZ0Z_23;
    wire un2_r_count_5hz_1_cry_22;
    wire r_count_5hzZ0Z_24;
    wire un2_r_count_5hz_1_cry_23;
    wire un2_r_count_5hz_1_cry_24;
    wire r_count_5hzZ0Z_25;
    wire bfn_9_5_0_;
    wire r_count_5hzZ0Z_26;
    wire un2_r_count_5hz_1_cry_25;
    wire r_count_5hzZ0Z_27;
    wire un2_r_count_5hz_1_cry_26;
    wire r_count_5hzZ0Z_28;
    wire un2_r_count_5hz_1_cry_27;
    wire r_count_5hzZ0Z_29;
    wire un2_r_count_5hz_1_cry_28;
    wire r_count_5hzZ0Z_30;
    wire un2_r_count_5hz_1_cry_29;
    wire un2_r_count_5hz_1_cry_30;
    wire r_count_5hzZ0Z_31;
    wire o_LED_43_0_and;
    wire bfn_9_9_0_;
    wire o_LED_43_0;
    wire o_LED_43_1;
    wire o_LED_43_3_and;
    wire o_LED_43_2;
    wire o_LED_43_3;
    wire o_LED_43_4;
    wire o_LED_43_5;
    wire o_LED_43_6;
    wire o_LED_43;
    wire bfn_9_10_0_;
    wire o_LED_43_THRU_CO_cascade_;
    wire o_LED_43_1_and;
    wire o_LED_43_2_and;
    wire o_LED_43_THRU_CO;
    wire bfn_11_1_0_;
    wire o_LED_13_0;
    wire o_LED_13_1;
    wire o_LED_13_2;
    wire o_LED_13_3;
    wire o_LED_13_4;
    wire o_LED_13_5;
    wire o_LED_13_6;
    wire o_LED_13;
    wire bfn_11_2_0_;
    wire o_LED_13_THRU_CO_cascade_;
    wire o_LED_13_1_and;
    wire o_LED_1_c;
    wire o_LED_13_4_and;
    wire o_LED_13_5_and;
    wire o_LED_13_6_and;
    wire o_LED_13_7_and;
    wire o_LED_43_4_and;
    wire r_count_1hzZ0Z_0;
    wire r_count_1hzZ0Z_1;
    wire bfn_11_9_0_;
    wire r_count_1hzZ0Z_2;
    wire un2_r_count_1hz_1_cry_1;
    wire r_count_1hzZ0Z_3;
    wire un2_r_count_1hz_1_cry_2;
    wire r_count_1hzZ0Z_4;
    wire un2_r_count_1hz_1_cry_3;
    wire r_count_1hzZ0Z_5;
    wire un2_r_count_1hz_1_cry_4_THRU_CO;
    wire un2_r_count_1hz_1_cry_4;
    wire r_count_1hzZ0Z_6;
    wire un2_r_count_1hz_1_cry_5;
    wire r_count_1hzZ0Z_7;
    wire un2_r_count_1hz_1_cry_6;
    wire r_count_1hzZ0Z_8;
    wire un2_r_count_1hz_1_cry_7;
    wire un2_r_count_1hz_1_cry_8;
    wire bfn_11_10_0_;
    wire r_count_1hzZ0Z_10;
    wire un2_r_count_1hz_1_cry_9_THRU_CO;
    wire un2_r_count_1hz_1_cry_9;
    wire r_count_1hzZ0Z_11;
    wire un2_r_count_1hz_1_cry_10_THRU_CO;
    wire un2_r_count_1hz_1_cry_10;
    wire r_count_1hzZ0Z_12;
    wire un2_r_count_1hz_1_cry_11_THRU_CO;
    wire un2_r_count_1hz_1_cry_11;
    wire r_count_1hzZ0Z_13;
    wire un2_r_count_1hz_1_cry_12_THRU_CO;
    wire un2_r_count_1hz_1_cry_12;
    wire un2_r_count_1hz_1_cry_13;
    wire r_count_1hzZ0Z_15;
    wire un2_r_count_1hz_1_cry_14_THRU_CO;
    wire un2_r_count_1hz_1_cry_14;
    wire un2_r_count_1hz_1_cry_15;
    wire un2_r_count_1hz_1_cry_16;
    wire r_count_1hzZ0Z_17;
    wire un2_r_count_1hz_1_cry_16_THRU_CO;
    wire bfn_11_11_0_;
    wire r_count_1hzZ0Z_18;
    wire un2_r_count_1hz_1_cry_17_THRU_CO;
    wire un2_r_count_1hz_1_cry_17;
    wire r_count_1hzZ0Z_19;
    wire un2_r_count_1hz_1_cry_18_THRU_CO;
    wire un2_r_count_1hz_1_cry_18;
    wire r_count_1hzZ0Z_20;
    wire un2_r_count_1hz_1_cry_19_THRU_CO;
    wire un2_r_count_1hz_1_cry_19;
    wire r_count_1hzZ0Z_21;
    wire un2_r_count_1hz_1_cry_20_THRU_CO;
    wire un2_r_count_1hz_1_cry_20;
    wire un2_r_count_1hz_1_cry_21;
    wire r_count_1hzZ0Z_23;
    wire un2_r_count_1hz_1_cry_22_THRU_CO;
    wire un2_r_count_1hz_1_cry_22;
    wire un2_r_count_1hz_1_cry_23;
    wire un2_r_count_1hz_1_cry_24;
    wire bfn_11_12_0_;
    wire un2_r_count_1hz_1_cry_25;
    wire un2_r_count_1hz_1_cry_26;
    wire un2_r_count_1hz_1_cry_27;
    wire un2_r_count_1hz_1_cry_28;
    wire un2_r_count_1hz_1_cry_29;
    wire un2_r_count_1hz_1_cry_30;
    wire r_count_1hzZ0Z_29;
    wire r_count_1hzZ0Z_31;
    wire r_count_1hzZ0Z_28;
    wire r_count_1hzZ0Z_30;
    wire o_LED_43_7_and;
    wire o_LED_13_THRU_CO;
    wire o_LED_13_0_and;
    wire o_LED_13_3_and;
    wire o_LED_13_2_and;
    wire r_count_10hzZ0Z_0;
    wire r_count_10hzZ0Z_1;
    wire bfn_12_3_0_;
    wire r_count_10hzZ0Z_2;
    wire un2_r_count_10hz_1_cry_1;
    wire r_count_10hzZ0Z_3;
    wire un2_r_count_10hz_1_cry_2;
    wire r_count_10hzZ0Z_4;
    wire un2_r_count_10hz_1_cry_3_THRU_CO;
    wire un2_r_count_10hz_1_cry_3;
    wire r_count_10hzZ0Z_5;
    wire un2_r_count_10hz_1_cry_4;
    wire r_count_10hzZ0Z_6;
    wire un2_r_count_10hz_1_cry_5_THRU_CO;
    wire un2_r_count_10hz_1_cry_5;
    wire r_count_10hzZ0Z_7;
    wire un2_r_count_10hz_1_cry_6_THRU_CO;
    wire un2_r_count_10hz_1_cry_6;
    wire r_count_10hzZ0Z_8;
    wire un2_r_count_10hz_1_cry_7;
    wire un2_r_count_10hz_1_cry_8;
    wire r_count_10hzZ0Z_9;
    wire un2_r_count_10hz_1_cry_8_THRU_CO;
    wire bfn_12_4_0_;
    wire r_count_10hzZ0Z_10;
    wire un2_r_count_10hz_1_cry_9;
    wire r_count_10hzZ0Z_11;
    wire un2_r_count_10hz_1_cry_10;
    wire r_count_10hzZ0Z_12;
    wire un2_r_count_10hz_1_cry_11_THRU_CO;
    wire un2_r_count_10hz_1_cry_11;
    wire r_count_10hzZ0Z_13;
    wire un2_r_count_10hz_1_cry_12;
    wire r_count_10hzZ0Z_14;
    wire un2_r_count_10hz_1_cry_13;
    wire r_count_10hzZ0Z_15;
    wire un2_r_count_10hz_1_cry_14;
    wire r_count_10hzZ0Z_16;
    wire un2_r_count_10hz_1_cry_15_THRU_CO;
    wire un2_r_count_10hz_1_cry_15;
    wire un2_r_count_10hz_1_cry_16;
    wire r_count_10hzZ0Z_17;
    wire un2_r_count_10hz_1_cry_16_THRU_CO;
    wire bfn_12_5_0_;
    wire r_count_10hzZ0Z_18;
    wire un2_r_count_10hz_1_cry_17;
    wire r_count_10hzZ0Z_19;
    wire un2_r_count_10hz_1_cry_18;
    wire r_count_10hzZ0Z_20;
    wire un2_r_count_10hz_1_cry_19_THRU_CO;
    wire un2_r_count_10hz_1_cry_19;
    wire r_count_10hzZ0Z_21;
    wire un2_r_count_10hz_1_cry_20;
    wire r_count_10hzZ0Z_22;
    wire un2_r_count_10hz_1_cry_21;
    wire r_count_10hzZ0Z_23;
    wire un2_r_count_10hz_1_cry_22;
    wire r_count_10hzZ0Z_24;
    wire un2_r_count_10hz_1_cry_23;
    wire un2_r_count_10hz_1_cry_24;
    wire r_count_10hzZ0Z_25;
    wire bfn_12_6_0_;
    wire r_count_10hzZ0Z_26;
    wire un2_r_count_10hz_1_cry_25;
    wire r_count_10hzZ0Z_27;
    wire un2_r_count_10hz_1_cry_26;
    wire r_count_10hzZ0Z_28;
    wire un2_r_count_10hz_1_cry_27;
    wire r_count_10hzZ0Z_29;
    wire un2_r_count_10hz_1_cry_28;
    wire r_count_10hzZ0Z_30;
    wire un2_r_count_10hz_1_cry_29;
    wire un2_r_count_10hz_1_cry_30;
    wire r_count_10hzZ0Z_31;
    wire i_Clk_c_g;
    wire r_count_1hzZ0Z_14;
    wire r_count_1hzZ0Z_22;
    wire r_count_1hzZ0Z_9;
    wire r_count_1hzZ0Z_16;
    wire o_LED_43_5_and;
    wire r_count_1hzZ0Z_25;
    wire r_count_1hzZ0Z_26;
    wire r_count_1hzZ0Z_24;
    wire r_count_1hzZ0Z_27;
    wire o_LED_43_6_and;
    wire _gnd_net_;

    PRE_IO_GBUF i_Clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__6647),
            .GLOBALBUFFEROUTPUT(i_Clk_c_g));
    IO_PAD i_Clk_ibuf_gb_io_iopad (
            .OE(N__6649),
            .DIN(N__6648),
            .DOUT(N__6647),
            .PACKAGEPIN(i_Clk));
    defparam i_Clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam i_Clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO i_Clk_ibuf_gb_io_preio (
            .PADOEN(N__6649),
            .PADOUT(N__6648),
            .PADIN(N__6647),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_1_obuf_iopad (
            .OE(N__6638),
            .DIN(N__6637),
            .DOUT(N__6636),
            .PACKAGEPIN(o_LED_1));
    defparam o_LED_1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_1_obuf_preio (
            .PADOEN(N__6638),
            .PADOUT(N__6637),
            .PADIN(N__6636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4954),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_2_obuf_iopad (
            .OE(N__6629),
            .DIN(N__6628),
            .DOUT(N__6627),
            .PACKAGEPIN(o_LED_2));
    defparam o_LED_2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_2_obuf_preio (
            .PADOEN(N__6629),
            .PADOUT(N__6628),
            .PADIN(N__6627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3376),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_4_obuf_iopad (
            .OE(N__6620),
            .DIN(N__6619),
            .DOUT(N__6618),
            .PACKAGEPIN(o_LED_4));
    defparam o_LED_4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_4_obuf_preio (
            .PADOEN(N__6620),
            .PADOUT(N__6619),
            .PADIN(N__6618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4228),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_LED_3_obuf_iopad (
            .OE(N__6611),
            .DIN(N__6610),
            .DOUT(N__6609),
            .PACKAGEPIN(o_LED_3));
    defparam o_LED_3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_LED_3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_LED_3_obuf_preio (
            .PADOEN(N__6611),
            .PADOUT(N__6610),
            .PADIN(N__6609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3208),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1415 (
            .O(N__6592),
            .I(N__6588));
    InMux I__1414 (
            .O(N__6591),
            .I(N__6585));
    LocalMux I__1413 (
            .O(N__6588),
            .I(r_count_10hzZ0Z_27));
    LocalMux I__1412 (
            .O(N__6585),
            .I(r_count_10hzZ0Z_27));
    InMux I__1411 (
            .O(N__6580),
            .I(un2_r_count_10hz_1_cry_26));
    CascadeMux I__1410 (
            .O(N__6577),
            .I(N__6573));
    InMux I__1409 (
            .O(N__6576),
            .I(N__6570));
    InMux I__1408 (
            .O(N__6573),
            .I(N__6567));
    LocalMux I__1407 (
            .O(N__6570),
            .I(r_count_10hzZ0Z_28));
    LocalMux I__1406 (
            .O(N__6567),
            .I(r_count_10hzZ0Z_28));
    InMux I__1405 (
            .O(N__6562),
            .I(un2_r_count_10hz_1_cry_27));
    InMux I__1404 (
            .O(N__6559),
            .I(N__6555));
    InMux I__1403 (
            .O(N__6558),
            .I(N__6552));
    LocalMux I__1402 (
            .O(N__6555),
            .I(r_count_10hzZ0Z_29));
    LocalMux I__1401 (
            .O(N__6552),
            .I(r_count_10hzZ0Z_29));
    InMux I__1400 (
            .O(N__6547),
            .I(un2_r_count_10hz_1_cry_28));
    InMux I__1399 (
            .O(N__6544),
            .I(N__6540));
    InMux I__1398 (
            .O(N__6543),
            .I(N__6537));
    LocalMux I__1397 (
            .O(N__6540),
            .I(r_count_10hzZ0Z_30));
    LocalMux I__1396 (
            .O(N__6537),
            .I(r_count_10hzZ0Z_30));
    InMux I__1395 (
            .O(N__6532),
            .I(un2_r_count_10hz_1_cry_29));
    InMux I__1394 (
            .O(N__6529),
            .I(un2_r_count_10hz_1_cry_30));
    InMux I__1393 (
            .O(N__6526),
            .I(N__6522));
    InMux I__1392 (
            .O(N__6525),
            .I(N__6519));
    LocalMux I__1391 (
            .O(N__6522),
            .I(r_count_10hzZ0Z_31));
    LocalMux I__1390 (
            .O(N__6519),
            .I(r_count_10hzZ0Z_31));
    ClkMux I__1389 (
            .O(N__6514),
            .I(N__6421));
    ClkMux I__1388 (
            .O(N__6513),
            .I(N__6421));
    ClkMux I__1387 (
            .O(N__6512),
            .I(N__6421));
    ClkMux I__1386 (
            .O(N__6511),
            .I(N__6421));
    ClkMux I__1385 (
            .O(N__6510),
            .I(N__6421));
    ClkMux I__1384 (
            .O(N__6509),
            .I(N__6421));
    ClkMux I__1383 (
            .O(N__6508),
            .I(N__6421));
    ClkMux I__1382 (
            .O(N__6507),
            .I(N__6421));
    ClkMux I__1381 (
            .O(N__6506),
            .I(N__6421));
    ClkMux I__1380 (
            .O(N__6505),
            .I(N__6421));
    ClkMux I__1379 (
            .O(N__6504),
            .I(N__6421));
    ClkMux I__1378 (
            .O(N__6503),
            .I(N__6421));
    ClkMux I__1377 (
            .O(N__6502),
            .I(N__6421));
    ClkMux I__1376 (
            .O(N__6501),
            .I(N__6421));
    ClkMux I__1375 (
            .O(N__6500),
            .I(N__6421));
    ClkMux I__1374 (
            .O(N__6499),
            .I(N__6421));
    ClkMux I__1373 (
            .O(N__6498),
            .I(N__6421));
    ClkMux I__1372 (
            .O(N__6497),
            .I(N__6421));
    ClkMux I__1371 (
            .O(N__6496),
            .I(N__6421));
    ClkMux I__1370 (
            .O(N__6495),
            .I(N__6421));
    ClkMux I__1369 (
            .O(N__6494),
            .I(N__6421));
    ClkMux I__1368 (
            .O(N__6493),
            .I(N__6421));
    ClkMux I__1367 (
            .O(N__6492),
            .I(N__6421));
    ClkMux I__1366 (
            .O(N__6491),
            .I(N__6421));
    ClkMux I__1365 (
            .O(N__6490),
            .I(N__6421));
    ClkMux I__1364 (
            .O(N__6489),
            .I(N__6421));
    ClkMux I__1363 (
            .O(N__6488),
            .I(N__6421));
    ClkMux I__1362 (
            .O(N__6487),
            .I(N__6421));
    ClkMux I__1361 (
            .O(N__6486),
            .I(N__6421));
    ClkMux I__1360 (
            .O(N__6485),
            .I(N__6421));
    ClkMux I__1359 (
            .O(N__6484),
            .I(N__6421));
    GlobalMux I__1358 (
            .O(N__6421),
            .I(N__6418));
    gio2CtrlBuf I__1357 (
            .O(N__6418),
            .I(i_Clk_c_g));
    InMux I__1356 (
            .O(N__6415),
            .I(N__6411));
    InMux I__1355 (
            .O(N__6414),
            .I(N__6408));
    LocalMux I__1354 (
            .O(N__6411),
            .I(r_count_1hzZ0Z_14));
    LocalMux I__1353 (
            .O(N__6408),
            .I(r_count_1hzZ0Z_14));
    InMux I__1352 (
            .O(N__6403),
            .I(N__6399));
    InMux I__1351 (
            .O(N__6402),
            .I(N__6396));
    LocalMux I__1350 (
            .O(N__6399),
            .I(r_count_1hzZ0Z_22));
    LocalMux I__1349 (
            .O(N__6396),
            .I(r_count_1hzZ0Z_22));
    CascadeMux I__1348 (
            .O(N__6391),
            .I(N__6387));
    InMux I__1347 (
            .O(N__6390),
            .I(N__6384));
    InMux I__1346 (
            .O(N__6387),
            .I(N__6381));
    LocalMux I__1345 (
            .O(N__6384),
            .I(r_count_1hzZ0Z_9));
    LocalMux I__1344 (
            .O(N__6381),
            .I(r_count_1hzZ0Z_9));
    InMux I__1343 (
            .O(N__6376),
            .I(N__6372));
    InMux I__1342 (
            .O(N__6375),
            .I(N__6369));
    LocalMux I__1341 (
            .O(N__6372),
            .I(r_count_1hzZ0Z_16));
    LocalMux I__1340 (
            .O(N__6369),
            .I(r_count_1hzZ0Z_16));
    InMux I__1339 (
            .O(N__6364),
            .I(N__6361));
    LocalMux I__1338 (
            .O(N__6361),
            .I(N__6358));
    Span4Mux_v I__1337 (
            .O(N__6358),
            .I(N__6355));
    Odrv4 I__1336 (
            .O(N__6355),
            .I(o_LED_43_5_and));
    InMux I__1335 (
            .O(N__6352),
            .I(N__6348));
    InMux I__1334 (
            .O(N__6351),
            .I(N__6345));
    LocalMux I__1333 (
            .O(N__6348),
            .I(r_count_1hzZ0Z_25));
    LocalMux I__1332 (
            .O(N__6345),
            .I(r_count_1hzZ0Z_25));
    InMux I__1331 (
            .O(N__6340),
            .I(N__6336));
    InMux I__1330 (
            .O(N__6339),
            .I(N__6333));
    LocalMux I__1329 (
            .O(N__6336),
            .I(r_count_1hzZ0Z_26));
    LocalMux I__1328 (
            .O(N__6333),
            .I(r_count_1hzZ0Z_26));
    CascadeMux I__1327 (
            .O(N__6328),
            .I(N__6324));
    InMux I__1326 (
            .O(N__6327),
            .I(N__6321));
    InMux I__1325 (
            .O(N__6324),
            .I(N__6318));
    LocalMux I__1324 (
            .O(N__6321),
            .I(r_count_1hzZ0Z_24));
    LocalMux I__1323 (
            .O(N__6318),
            .I(r_count_1hzZ0Z_24));
    InMux I__1322 (
            .O(N__6313),
            .I(N__6309));
    InMux I__1321 (
            .O(N__6312),
            .I(N__6306));
    LocalMux I__1320 (
            .O(N__6309),
            .I(r_count_1hzZ0Z_27));
    LocalMux I__1319 (
            .O(N__6306),
            .I(r_count_1hzZ0Z_27));
    CascadeMux I__1318 (
            .O(N__6301),
            .I(N__6298));
    InMux I__1317 (
            .O(N__6298),
            .I(N__6295));
    LocalMux I__1316 (
            .O(N__6295),
            .I(N__6292));
    Span4Mux_v I__1315 (
            .O(N__6292),
            .I(N__6289));
    Odrv4 I__1314 (
            .O(N__6289),
            .I(o_LED_43_6_and));
    InMux I__1313 (
            .O(N__6286),
            .I(N__6282));
    InMux I__1312 (
            .O(N__6285),
            .I(N__6279));
    LocalMux I__1311 (
            .O(N__6282),
            .I(N__6274));
    LocalMux I__1310 (
            .O(N__6279),
            .I(N__6274));
    Odrv4 I__1309 (
            .O(N__6274),
            .I(r_count_10hzZ0Z_19));
    InMux I__1308 (
            .O(N__6271),
            .I(un2_r_count_10hz_1_cry_18));
    InMux I__1307 (
            .O(N__6268),
            .I(N__6264));
    InMux I__1306 (
            .O(N__6267),
            .I(N__6260));
    LocalMux I__1305 (
            .O(N__6264),
            .I(N__6257));
    InMux I__1304 (
            .O(N__6263),
            .I(N__6254));
    LocalMux I__1303 (
            .O(N__6260),
            .I(r_count_10hzZ0Z_20));
    Odrv4 I__1302 (
            .O(N__6257),
            .I(r_count_10hzZ0Z_20));
    LocalMux I__1301 (
            .O(N__6254),
            .I(r_count_10hzZ0Z_20));
    InMux I__1300 (
            .O(N__6247),
            .I(N__6244));
    LocalMux I__1299 (
            .O(N__6244),
            .I(N__6241));
    Odrv4 I__1298 (
            .O(N__6241),
            .I(un2_r_count_10hz_1_cry_19_THRU_CO));
    InMux I__1297 (
            .O(N__6238),
            .I(un2_r_count_10hz_1_cry_19));
    InMux I__1296 (
            .O(N__6235),
            .I(N__6231));
    InMux I__1295 (
            .O(N__6234),
            .I(N__6228));
    LocalMux I__1294 (
            .O(N__6231),
            .I(N__6225));
    LocalMux I__1293 (
            .O(N__6228),
            .I(r_count_10hzZ0Z_21));
    Odrv4 I__1292 (
            .O(N__6225),
            .I(r_count_10hzZ0Z_21));
    InMux I__1291 (
            .O(N__6220),
            .I(un2_r_count_10hz_1_cry_20));
    CascadeMux I__1290 (
            .O(N__6217),
            .I(N__6214));
    InMux I__1289 (
            .O(N__6214),
            .I(N__6210));
    InMux I__1288 (
            .O(N__6213),
            .I(N__6207));
    LocalMux I__1287 (
            .O(N__6210),
            .I(N__6204));
    LocalMux I__1286 (
            .O(N__6207),
            .I(r_count_10hzZ0Z_22));
    Odrv4 I__1285 (
            .O(N__6204),
            .I(r_count_10hzZ0Z_22));
    InMux I__1284 (
            .O(N__6199),
            .I(un2_r_count_10hz_1_cry_21));
    InMux I__1283 (
            .O(N__6196),
            .I(N__6192));
    InMux I__1282 (
            .O(N__6195),
            .I(N__6189));
    LocalMux I__1281 (
            .O(N__6192),
            .I(r_count_10hzZ0Z_23));
    LocalMux I__1280 (
            .O(N__6189),
            .I(r_count_10hzZ0Z_23));
    InMux I__1279 (
            .O(N__6184),
            .I(un2_r_count_10hz_1_cry_22));
    InMux I__1278 (
            .O(N__6181),
            .I(N__6177));
    InMux I__1277 (
            .O(N__6180),
            .I(N__6174));
    LocalMux I__1276 (
            .O(N__6177),
            .I(r_count_10hzZ0Z_24));
    LocalMux I__1275 (
            .O(N__6174),
            .I(r_count_10hzZ0Z_24));
    InMux I__1274 (
            .O(N__6169),
            .I(un2_r_count_10hz_1_cry_23));
    CascadeMux I__1273 (
            .O(N__6166),
            .I(N__6162));
    InMux I__1272 (
            .O(N__6165),
            .I(N__6159));
    InMux I__1271 (
            .O(N__6162),
            .I(N__6156));
    LocalMux I__1270 (
            .O(N__6159),
            .I(r_count_10hzZ0Z_25));
    LocalMux I__1269 (
            .O(N__6156),
            .I(r_count_10hzZ0Z_25));
    InMux I__1268 (
            .O(N__6151),
            .I(bfn_12_6_0_));
    InMux I__1267 (
            .O(N__6148),
            .I(N__6144));
    InMux I__1266 (
            .O(N__6147),
            .I(N__6141));
    LocalMux I__1265 (
            .O(N__6144),
            .I(r_count_10hzZ0Z_26));
    LocalMux I__1264 (
            .O(N__6141),
            .I(r_count_10hzZ0Z_26));
    InMux I__1263 (
            .O(N__6136),
            .I(un2_r_count_10hz_1_cry_25));
    InMux I__1262 (
            .O(N__6133),
            .I(un2_r_count_10hz_1_cry_9));
    InMux I__1261 (
            .O(N__6130),
            .I(N__6126));
    InMux I__1260 (
            .O(N__6129),
            .I(N__6123));
    LocalMux I__1259 (
            .O(N__6126),
            .I(N__6120));
    LocalMux I__1258 (
            .O(N__6123),
            .I(r_count_10hzZ0Z_11));
    Odrv4 I__1257 (
            .O(N__6120),
            .I(r_count_10hzZ0Z_11));
    InMux I__1256 (
            .O(N__6115),
            .I(un2_r_count_10hz_1_cry_10));
    CascadeMux I__1255 (
            .O(N__6112),
            .I(N__6107));
    InMux I__1254 (
            .O(N__6111),
            .I(N__6104));
    InMux I__1253 (
            .O(N__6110),
            .I(N__6101));
    InMux I__1252 (
            .O(N__6107),
            .I(N__6098));
    LocalMux I__1251 (
            .O(N__6104),
            .I(r_count_10hzZ0Z_12));
    LocalMux I__1250 (
            .O(N__6101),
            .I(r_count_10hzZ0Z_12));
    LocalMux I__1249 (
            .O(N__6098),
            .I(r_count_10hzZ0Z_12));
    InMux I__1248 (
            .O(N__6091),
            .I(N__6088));
    LocalMux I__1247 (
            .O(N__6088),
            .I(un2_r_count_10hz_1_cry_11_THRU_CO));
    InMux I__1246 (
            .O(N__6085),
            .I(un2_r_count_10hz_1_cry_11));
    InMux I__1245 (
            .O(N__6082),
            .I(N__6078));
    InMux I__1244 (
            .O(N__6081),
            .I(N__6075));
    LocalMux I__1243 (
            .O(N__6078),
            .I(r_count_10hzZ0Z_13));
    LocalMux I__1242 (
            .O(N__6075),
            .I(r_count_10hzZ0Z_13));
    InMux I__1241 (
            .O(N__6070),
            .I(un2_r_count_10hz_1_cry_12));
    InMux I__1240 (
            .O(N__6067),
            .I(N__6063));
    InMux I__1239 (
            .O(N__6066),
            .I(N__6060));
    LocalMux I__1238 (
            .O(N__6063),
            .I(r_count_10hzZ0Z_14));
    LocalMux I__1237 (
            .O(N__6060),
            .I(r_count_10hzZ0Z_14));
    InMux I__1236 (
            .O(N__6055),
            .I(un2_r_count_10hz_1_cry_13));
    InMux I__1235 (
            .O(N__6052),
            .I(N__6048));
    InMux I__1234 (
            .O(N__6051),
            .I(N__6045));
    LocalMux I__1233 (
            .O(N__6048),
            .I(r_count_10hzZ0Z_15));
    LocalMux I__1232 (
            .O(N__6045),
            .I(r_count_10hzZ0Z_15));
    InMux I__1231 (
            .O(N__6040),
            .I(un2_r_count_10hz_1_cry_14));
    InMux I__1230 (
            .O(N__6037),
            .I(N__6032));
    InMux I__1229 (
            .O(N__6036),
            .I(N__6029));
    InMux I__1228 (
            .O(N__6035),
            .I(N__6026));
    LocalMux I__1227 (
            .O(N__6032),
            .I(r_count_10hzZ0Z_16));
    LocalMux I__1226 (
            .O(N__6029),
            .I(r_count_10hzZ0Z_16));
    LocalMux I__1225 (
            .O(N__6026),
            .I(r_count_10hzZ0Z_16));
    InMux I__1224 (
            .O(N__6019),
            .I(N__6016));
    LocalMux I__1223 (
            .O(N__6016),
            .I(un2_r_count_10hz_1_cry_15_THRU_CO));
    InMux I__1222 (
            .O(N__6013),
            .I(un2_r_count_10hz_1_cry_15));
    InMux I__1221 (
            .O(N__6010),
            .I(N__6006));
    InMux I__1220 (
            .O(N__6009),
            .I(N__6002));
    LocalMux I__1219 (
            .O(N__6006),
            .I(N__5999));
    InMux I__1218 (
            .O(N__6005),
            .I(N__5996));
    LocalMux I__1217 (
            .O(N__6002),
            .I(r_count_10hzZ0Z_17));
    Odrv4 I__1216 (
            .O(N__5999),
            .I(r_count_10hzZ0Z_17));
    LocalMux I__1215 (
            .O(N__5996),
            .I(r_count_10hzZ0Z_17));
    InMux I__1214 (
            .O(N__5989),
            .I(N__5986));
    LocalMux I__1213 (
            .O(N__5986),
            .I(N__5983));
    Odrv4 I__1212 (
            .O(N__5983),
            .I(un2_r_count_10hz_1_cry_16_THRU_CO));
    InMux I__1211 (
            .O(N__5980),
            .I(bfn_12_5_0_));
    CascadeMux I__1210 (
            .O(N__5977),
            .I(N__5973));
    InMux I__1209 (
            .O(N__5976),
            .I(N__5970));
    InMux I__1208 (
            .O(N__5973),
            .I(N__5967));
    LocalMux I__1207 (
            .O(N__5970),
            .I(r_count_10hzZ0Z_18));
    LocalMux I__1206 (
            .O(N__5967),
            .I(r_count_10hzZ0Z_18));
    InMux I__1205 (
            .O(N__5962),
            .I(un2_r_count_10hz_1_cry_17));
    InMux I__1204 (
            .O(N__5959),
            .I(N__5955));
    InMux I__1203 (
            .O(N__5958),
            .I(N__5952));
    LocalMux I__1202 (
            .O(N__5955),
            .I(r_count_10hzZ0Z_2));
    LocalMux I__1201 (
            .O(N__5952),
            .I(r_count_10hzZ0Z_2));
    InMux I__1200 (
            .O(N__5947),
            .I(un2_r_count_10hz_1_cry_1));
    InMux I__1199 (
            .O(N__5944),
            .I(N__5940));
    InMux I__1198 (
            .O(N__5943),
            .I(N__5937));
    LocalMux I__1197 (
            .O(N__5940),
            .I(r_count_10hzZ0Z_3));
    LocalMux I__1196 (
            .O(N__5937),
            .I(r_count_10hzZ0Z_3));
    InMux I__1195 (
            .O(N__5932),
            .I(un2_r_count_10hz_1_cry_2));
    InMux I__1194 (
            .O(N__5929),
            .I(N__5924));
    InMux I__1193 (
            .O(N__5928),
            .I(N__5921));
    InMux I__1192 (
            .O(N__5927),
            .I(N__5918));
    LocalMux I__1191 (
            .O(N__5924),
            .I(r_count_10hzZ0Z_4));
    LocalMux I__1190 (
            .O(N__5921),
            .I(r_count_10hzZ0Z_4));
    LocalMux I__1189 (
            .O(N__5918),
            .I(r_count_10hzZ0Z_4));
    InMux I__1188 (
            .O(N__5911),
            .I(N__5908));
    LocalMux I__1187 (
            .O(N__5908),
            .I(un2_r_count_10hz_1_cry_3_THRU_CO));
    InMux I__1186 (
            .O(N__5905),
            .I(un2_r_count_10hz_1_cry_3));
    InMux I__1185 (
            .O(N__5902),
            .I(N__5898));
    InMux I__1184 (
            .O(N__5901),
            .I(N__5895));
    LocalMux I__1183 (
            .O(N__5898),
            .I(r_count_10hzZ0Z_5));
    LocalMux I__1182 (
            .O(N__5895),
            .I(r_count_10hzZ0Z_5));
    InMux I__1181 (
            .O(N__5890),
            .I(un2_r_count_10hz_1_cry_4));
    InMux I__1180 (
            .O(N__5887),
            .I(N__5882));
    InMux I__1179 (
            .O(N__5886),
            .I(N__5879));
    InMux I__1178 (
            .O(N__5885),
            .I(N__5876));
    LocalMux I__1177 (
            .O(N__5882),
            .I(r_count_10hzZ0Z_6));
    LocalMux I__1176 (
            .O(N__5879),
            .I(r_count_10hzZ0Z_6));
    LocalMux I__1175 (
            .O(N__5876),
            .I(r_count_10hzZ0Z_6));
    InMux I__1174 (
            .O(N__5869),
            .I(N__5866));
    LocalMux I__1173 (
            .O(N__5866),
            .I(un2_r_count_10hz_1_cry_5_THRU_CO));
    InMux I__1172 (
            .O(N__5863),
            .I(un2_r_count_10hz_1_cry_5));
    CascadeMux I__1171 (
            .O(N__5860),
            .I(N__5856));
    InMux I__1170 (
            .O(N__5859),
            .I(N__5850));
    InMux I__1169 (
            .O(N__5856),
            .I(N__5850));
    InMux I__1168 (
            .O(N__5855),
            .I(N__5847));
    LocalMux I__1167 (
            .O(N__5850),
            .I(r_count_10hzZ0Z_7));
    LocalMux I__1166 (
            .O(N__5847),
            .I(r_count_10hzZ0Z_7));
    InMux I__1165 (
            .O(N__5842),
            .I(N__5839));
    LocalMux I__1164 (
            .O(N__5839),
            .I(un2_r_count_10hz_1_cry_6_THRU_CO));
    InMux I__1163 (
            .O(N__5836),
            .I(un2_r_count_10hz_1_cry_6));
    InMux I__1162 (
            .O(N__5833),
            .I(N__5829));
    InMux I__1161 (
            .O(N__5832),
            .I(N__5826));
    LocalMux I__1160 (
            .O(N__5829),
            .I(r_count_10hzZ0Z_8));
    LocalMux I__1159 (
            .O(N__5826),
            .I(r_count_10hzZ0Z_8));
    InMux I__1158 (
            .O(N__5821),
            .I(un2_r_count_10hz_1_cry_7));
    InMux I__1157 (
            .O(N__5818),
            .I(N__5813));
    InMux I__1156 (
            .O(N__5817),
            .I(N__5810));
    InMux I__1155 (
            .O(N__5816),
            .I(N__5807));
    LocalMux I__1154 (
            .O(N__5813),
            .I(r_count_10hzZ0Z_9));
    LocalMux I__1153 (
            .O(N__5810),
            .I(r_count_10hzZ0Z_9));
    LocalMux I__1152 (
            .O(N__5807),
            .I(r_count_10hzZ0Z_9));
    InMux I__1151 (
            .O(N__5800),
            .I(N__5797));
    LocalMux I__1150 (
            .O(N__5797),
            .I(un2_r_count_10hz_1_cry_8_THRU_CO));
    InMux I__1149 (
            .O(N__5794),
            .I(bfn_12_4_0_));
    CascadeMux I__1148 (
            .O(N__5791),
            .I(N__5788));
    InMux I__1147 (
            .O(N__5788),
            .I(N__5784));
    InMux I__1146 (
            .O(N__5787),
            .I(N__5781));
    LocalMux I__1145 (
            .O(N__5784),
            .I(N__5778));
    LocalMux I__1144 (
            .O(N__5781),
            .I(r_count_10hzZ0Z_10));
    Odrv12 I__1143 (
            .O(N__5778),
            .I(r_count_10hzZ0Z_10));
    InMux I__1142 (
            .O(N__5773),
            .I(N__5767));
    InMux I__1141 (
            .O(N__5772),
            .I(N__5767));
    LocalMux I__1140 (
            .O(N__5767),
            .I(r_count_1hzZ0Z_31));
    CascadeMux I__1139 (
            .O(N__5764),
            .I(N__5760));
    CascadeMux I__1138 (
            .O(N__5763),
            .I(N__5757));
    InMux I__1137 (
            .O(N__5760),
            .I(N__5752));
    InMux I__1136 (
            .O(N__5757),
            .I(N__5752));
    LocalMux I__1135 (
            .O(N__5752),
            .I(r_count_1hzZ0Z_28));
    InMux I__1134 (
            .O(N__5749),
            .I(N__5743));
    InMux I__1133 (
            .O(N__5748),
            .I(N__5743));
    LocalMux I__1132 (
            .O(N__5743),
            .I(r_count_1hzZ0Z_30));
    CascadeMux I__1131 (
            .O(N__5740),
            .I(N__5737));
    InMux I__1130 (
            .O(N__5737),
            .I(N__5734));
    LocalMux I__1129 (
            .O(N__5734),
            .I(N__5731));
    Span4Mux_h I__1128 (
            .O(N__5731),
            .I(N__5728));
    Odrv4 I__1127 (
            .O(N__5728),
            .I(o_LED_43_7_and));
    CascadeMux I__1126 (
            .O(N__5725),
            .I(N__5717));
    CascadeMux I__1125 (
            .O(N__5724),
            .I(N__5711));
    CascadeMux I__1124 (
            .O(N__5723),
            .I(N__5708));
    CascadeMux I__1123 (
            .O(N__5722),
            .I(N__5705));
    CascadeMux I__1122 (
            .O(N__5721),
            .I(N__5702));
    InMux I__1121 (
            .O(N__5720),
            .I(N__5695));
    InMux I__1120 (
            .O(N__5717),
            .I(N__5695));
    InMux I__1119 (
            .O(N__5716),
            .I(N__5695));
    InMux I__1118 (
            .O(N__5715),
            .I(N__5682));
    InMux I__1117 (
            .O(N__5714),
            .I(N__5682));
    InMux I__1116 (
            .O(N__5711),
            .I(N__5682));
    InMux I__1115 (
            .O(N__5708),
            .I(N__5682));
    InMux I__1114 (
            .O(N__5705),
            .I(N__5682));
    InMux I__1113 (
            .O(N__5702),
            .I(N__5682));
    LocalMux I__1112 (
            .O(N__5695),
            .I(o_LED_13_THRU_CO));
    LocalMux I__1111 (
            .O(N__5682),
            .I(o_LED_13_THRU_CO));
    CascadeMux I__1110 (
            .O(N__5677),
            .I(N__5674));
    InMux I__1109 (
            .O(N__5674),
            .I(N__5671));
    LocalMux I__1108 (
            .O(N__5671),
            .I(o_LED_13_0_and));
    CascadeMux I__1107 (
            .O(N__5668),
            .I(N__5665));
    InMux I__1106 (
            .O(N__5665),
            .I(N__5662));
    LocalMux I__1105 (
            .O(N__5662),
            .I(o_LED_13_3_and));
    InMux I__1104 (
            .O(N__5659),
            .I(N__5656));
    LocalMux I__1103 (
            .O(N__5656),
            .I(o_LED_13_2_and));
    CascadeMux I__1102 (
            .O(N__5653),
            .I(N__5649));
    CascadeMux I__1101 (
            .O(N__5652),
            .I(N__5645));
    InMux I__1100 (
            .O(N__5649),
            .I(N__5637));
    InMux I__1099 (
            .O(N__5648),
            .I(N__5637));
    InMux I__1098 (
            .O(N__5645),
            .I(N__5637));
    InMux I__1097 (
            .O(N__5644),
            .I(N__5634));
    LocalMux I__1096 (
            .O(N__5637),
            .I(r_count_10hzZ0Z_0));
    LocalMux I__1095 (
            .O(N__5634),
            .I(r_count_10hzZ0Z_0));
    InMux I__1094 (
            .O(N__5629),
            .I(N__5622));
    InMux I__1093 (
            .O(N__5628),
            .I(N__5622));
    CascadeMux I__1092 (
            .O(N__5627),
            .I(N__5619));
    LocalMux I__1091 (
            .O(N__5622),
            .I(N__5616));
    InMux I__1090 (
            .O(N__5619),
            .I(N__5613));
    Odrv4 I__1089 (
            .O(N__5616),
            .I(r_count_10hzZ0Z_1));
    LocalMux I__1088 (
            .O(N__5613),
            .I(r_count_10hzZ0Z_1));
    InMux I__1087 (
            .O(N__5608),
            .I(un2_r_count_1hz_1_cry_22));
    InMux I__1086 (
            .O(N__5605),
            .I(un2_r_count_1hz_1_cry_23));
    InMux I__1085 (
            .O(N__5602),
            .I(bfn_11_12_0_));
    InMux I__1084 (
            .O(N__5599),
            .I(un2_r_count_1hz_1_cry_25));
    InMux I__1083 (
            .O(N__5596),
            .I(un2_r_count_1hz_1_cry_26));
    InMux I__1082 (
            .O(N__5593),
            .I(un2_r_count_1hz_1_cry_27));
    InMux I__1081 (
            .O(N__5590),
            .I(un2_r_count_1hz_1_cry_28));
    InMux I__1080 (
            .O(N__5587),
            .I(un2_r_count_1hz_1_cry_29));
    InMux I__1079 (
            .O(N__5584),
            .I(un2_r_count_1hz_1_cry_30));
    InMux I__1078 (
            .O(N__5581),
            .I(N__5575));
    InMux I__1077 (
            .O(N__5580),
            .I(N__5575));
    LocalMux I__1076 (
            .O(N__5575),
            .I(r_count_1hzZ0Z_29));
    InMux I__1075 (
            .O(N__5572),
            .I(N__5569));
    LocalMux I__1074 (
            .O(N__5569),
            .I(N__5566));
    Odrv4 I__1073 (
            .O(N__5566),
            .I(un2_r_count_1hz_1_cry_14_THRU_CO));
    InMux I__1072 (
            .O(N__5563),
            .I(un2_r_count_1hz_1_cry_14));
    InMux I__1071 (
            .O(N__5560),
            .I(un2_r_count_1hz_1_cry_15));
    InMux I__1070 (
            .O(N__5557),
            .I(N__5552));
    CascadeMux I__1069 (
            .O(N__5556),
            .I(N__5549));
    InMux I__1068 (
            .O(N__5555),
            .I(N__5546));
    LocalMux I__1067 (
            .O(N__5552),
            .I(N__5543));
    InMux I__1066 (
            .O(N__5549),
            .I(N__5540));
    LocalMux I__1065 (
            .O(N__5546),
            .I(r_count_1hzZ0Z_17));
    Odrv4 I__1064 (
            .O(N__5543),
            .I(r_count_1hzZ0Z_17));
    LocalMux I__1063 (
            .O(N__5540),
            .I(r_count_1hzZ0Z_17));
    InMux I__1062 (
            .O(N__5533),
            .I(N__5530));
    LocalMux I__1061 (
            .O(N__5530),
            .I(N__5527));
    Span4Mux_h I__1060 (
            .O(N__5527),
            .I(N__5524));
    Odrv4 I__1059 (
            .O(N__5524),
            .I(un2_r_count_1hz_1_cry_16_THRU_CO));
    InMux I__1058 (
            .O(N__5521),
            .I(bfn_11_11_0_));
    InMux I__1057 (
            .O(N__5518),
            .I(N__5514));
    InMux I__1056 (
            .O(N__5517),
            .I(N__5511));
    LocalMux I__1055 (
            .O(N__5514),
            .I(N__5505));
    LocalMux I__1054 (
            .O(N__5511),
            .I(N__5505));
    InMux I__1053 (
            .O(N__5510),
            .I(N__5502));
    Odrv4 I__1052 (
            .O(N__5505),
            .I(r_count_1hzZ0Z_18));
    LocalMux I__1051 (
            .O(N__5502),
            .I(r_count_1hzZ0Z_18));
    InMux I__1050 (
            .O(N__5497),
            .I(N__5494));
    LocalMux I__1049 (
            .O(N__5494),
            .I(N__5491));
    Span4Mux_h I__1048 (
            .O(N__5491),
            .I(N__5488));
    Odrv4 I__1047 (
            .O(N__5488),
            .I(un2_r_count_1hz_1_cry_17_THRU_CO));
    InMux I__1046 (
            .O(N__5485),
            .I(un2_r_count_1hz_1_cry_17));
    InMux I__1045 (
            .O(N__5482),
            .I(N__5478));
    InMux I__1044 (
            .O(N__5481),
            .I(N__5474));
    LocalMux I__1043 (
            .O(N__5478),
            .I(N__5471));
    InMux I__1042 (
            .O(N__5477),
            .I(N__5468));
    LocalMux I__1041 (
            .O(N__5474),
            .I(r_count_1hzZ0Z_19));
    Odrv4 I__1040 (
            .O(N__5471),
            .I(r_count_1hzZ0Z_19));
    LocalMux I__1039 (
            .O(N__5468),
            .I(r_count_1hzZ0Z_19));
    InMux I__1038 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__1037 (
            .O(N__5458),
            .I(N__5455));
    Span4Mux_h I__1036 (
            .O(N__5455),
            .I(N__5452));
    Odrv4 I__1035 (
            .O(N__5452),
            .I(un2_r_count_1hz_1_cry_18_THRU_CO));
    InMux I__1034 (
            .O(N__5449),
            .I(un2_r_count_1hz_1_cry_18));
    InMux I__1033 (
            .O(N__5446),
            .I(N__5442));
    InMux I__1032 (
            .O(N__5445),
            .I(N__5438));
    LocalMux I__1031 (
            .O(N__5442),
            .I(N__5435));
    InMux I__1030 (
            .O(N__5441),
            .I(N__5432));
    LocalMux I__1029 (
            .O(N__5438),
            .I(r_count_1hzZ0Z_20));
    Odrv4 I__1028 (
            .O(N__5435),
            .I(r_count_1hzZ0Z_20));
    LocalMux I__1027 (
            .O(N__5432),
            .I(r_count_1hzZ0Z_20));
    InMux I__1026 (
            .O(N__5425),
            .I(N__5422));
    LocalMux I__1025 (
            .O(N__5422),
            .I(N__5419));
    Odrv4 I__1024 (
            .O(N__5419),
            .I(un2_r_count_1hz_1_cry_19_THRU_CO));
    InMux I__1023 (
            .O(N__5416),
            .I(un2_r_count_1hz_1_cry_19));
    InMux I__1022 (
            .O(N__5413),
            .I(N__5408));
    CascadeMux I__1021 (
            .O(N__5412),
            .I(N__5405));
    InMux I__1020 (
            .O(N__5411),
            .I(N__5402));
    LocalMux I__1019 (
            .O(N__5408),
            .I(N__5399));
    InMux I__1018 (
            .O(N__5405),
            .I(N__5396));
    LocalMux I__1017 (
            .O(N__5402),
            .I(r_count_1hzZ0Z_21));
    Odrv12 I__1016 (
            .O(N__5399),
            .I(r_count_1hzZ0Z_21));
    LocalMux I__1015 (
            .O(N__5396),
            .I(r_count_1hzZ0Z_21));
    InMux I__1014 (
            .O(N__5389),
            .I(N__5386));
    LocalMux I__1013 (
            .O(N__5386),
            .I(N__5383));
    Odrv4 I__1012 (
            .O(N__5383),
            .I(un2_r_count_1hz_1_cry_20_THRU_CO));
    InMux I__1011 (
            .O(N__5380),
            .I(un2_r_count_1hz_1_cry_20));
    InMux I__1010 (
            .O(N__5377),
            .I(un2_r_count_1hz_1_cry_21));
    InMux I__1009 (
            .O(N__5374),
            .I(N__5369));
    InMux I__1008 (
            .O(N__5373),
            .I(N__5366));
    InMux I__1007 (
            .O(N__5372),
            .I(N__5363));
    LocalMux I__1006 (
            .O(N__5369),
            .I(N__5360));
    LocalMux I__1005 (
            .O(N__5366),
            .I(N__5357));
    LocalMux I__1004 (
            .O(N__5363),
            .I(r_count_1hzZ0Z_23));
    Odrv4 I__1003 (
            .O(N__5360),
            .I(r_count_1hzZ0Z_23));
    Odrv4 I__1002 (
            .O(N__5357),
            .I(r_count_1hzZ0Z_23));
    InMux I__1001 (
            .O(N__5350),
            .I(N__5347));
    LocalMux I__1000 (
            .O(N__5347),
            .I(N__5344));
    Odrv4 I__999 (
            .O(N__5344),
            .I(un2_r_count_1hz_1_cry_22_THRU_CO));
    CascadeMux I__998 (
            .O(N__5341),
            .I(N__5338));
    InMux I__997 (
            .O(N__5338),
            .I(N__5334));
    InMux I__996 (
            .O(N__5337),
            .I(N__5331));
    LocalMux I__995 (
            .O(N__5334),
            .I(r_count_1hzZ0Z_7));
    LocalMux I__994 (
            .O(N__5331),
            .I(r_count_1hzZ0Z_7));
    InMux I__993 (
            .O(N__5326),
            .I(un2_r_count_1hz_1_cry_6));
    InMux I__992 (
            .O(N__5323),
            .I(N__5319));
    InMux I__991 (
            .O(N__5322),
            .I(N__5316));
    LocalMux I__990 (
            .O(N__5319),
            .I(r_count_1hzZ0Z_8));
    LocalMux I__989 (
            .O(N__5316),
            .I(r_count_1hzZ0Z_8));
    InMux I__988 (
            .O(N__5311),
            .I(un2_r_count_1hz_1_cry_7));
    InMux I__987 (
            .O(N__5308),
            .I(bfn_11_10_0_));
    InMux I__986 (
            .O(N__5305),
            .I(N__5300));
    InMux I__985 (
            .O(N__5304),
            .I(N__5297));
    InMux I__984 (
            .O(N__5303),
            .I(N__5294));
    LocalMux I__983 (
            .O(N__5300),
            .I(N__5289));
    LocalMux I__982 (
            .O(N__5297),
            .I(N__5289));
    LocalMux I__981 (
            .O(N__5294),
            .I(r_count_1hzZ0Z_10));
    Odrv4 I__980 (
            .O(N__5289),
            .I(r_count_1hzZ0Z_10));
    InMux I__979 (
            .O(N__5284),
            .I(N__5281));
    LocalMux I__978 (
            .O(N__5281),
            .I(N__5278));
    Span4Mux_h I__977 (
            .O(N__5278),
            .I(N__5275));
    Odrv4 I__976 (
            .O(N__5275),
            .I(un2_r_count_1hz_1_cry_9_THRU_CO));
    InMux I__975 (
            .O(N__5272),
            .I(un2_r_count_1hz_1_cry_9));
    CascadeMux I__974 (
            .O(N__5269),
            .I(N__5264));
    InMux I__973 (
            .O(N__5268),
            .I(N__5261));
    InMux I__972 (
            .O(N__5267),
            .I(N__5258));
    InMux I__971 (
            .O(N__5264),
            .I(N__5255));
    LocalMux I__970 (
            .O(N__5261),
            .I(N__5252));
    LocalMux I__969 (
            .O(N__5258),
            .I(r_count_1hzZ0Z_11));
    LocalMux I__968 (
            .O(N__5255),
            .I(r_count_1hzZ0Z_11));
    Odrv4 I__967 (
            .O(N__5252),
            .I(r_count_1hzZ0Z_11));
    InMux I__966 (
            .O(N__5245),
            .I(N__5242));
    LocalMux I__965 (
            .O(N__5242),
            .I(N__5239));
    Span4Mux_h I__964 (
            .O(N__5239),
            .I(N__5236));
    Odrv4 I__963 (
            .O(N__5236),
            .I(un2_r_count_1hz_1_cry_10_THRU_CO));
    InMux I__962 (
            .O(N__5233),
            .I(un2_r_count_1hz_1_cry_10));
    InMux I__961 (
            .O(N__5230),
            .I(N__5226));
    InMux I__960 (
            .O(N__5229),
            .I(N__5222));
    LocalMux I__959 (
            .O(N__5226),
            .I(N__5219));
    InMux I__958 (
            .O(N__5225),
            .I(N__5216));
    LocalMux I__957 (
            .O(N__5222),
            .I(r_count_1hzZ0Z_12));
    Odrv4 I__956 (
            .O(N__5219),
            .I(r_count_1hzZ0Z_12));
    LocalMux I__955 (
            .O(N__5216),
            .I(r_count_1hzZ0Z_12));
    InMux I__954 (
            .O(N__5209),
            .I(N__5206));
    LocalMux I__953 (
            .O(N__5206),
            .I(N__5203));
    Span4Mux_h I__952 (
            .O(N__5203),
            .I(N__5200));
    Odrv4 I__951 (
            .O(N__5200),
            .I(un2_r_count_1hz_1_cry_11_THRU_CO));
    InMux I__950 (
            .O(N__5197),
            .I(un2_r_count_1hz_1_cry_11));
    InMux I__949 (
            .O(N__5194),
            .I(N__5189));
    InMux I__948 (
            .O(N__5193),
            .I(N__5184));
    InMux I__947 (
            .O(N__5192),
            .I(N__5184));
    LocalMux I__946 (
            .O(N__5189),
            .I(N__5181));
    LocalMux I__945 (
            .O(N__5184),
            .I(r_count_1hzZ0Z_13));
    Odrv4 I__944 (
            .O(N__5181),
            .I(r_count_1hzZ0Z_13));
    InMux I__943 (
            .O(N__5176),
            .I(N__5173));
    LocalMux I__942 (
            .O(N__5173),
            .I(N__5170));
    Odrv4 I__941 (
            .O(N__5170),
            .I(un2_r_count_1hz_1_cry_12_THRU_CO));
    InMux I__940 (
            .O(N__5167),
            .I(un2_r_count_1hz_1_cry_12));
    InMux I__939 (
            .O(N__5164),
            .I(un2_r_count_1hz_1_cry_13));
    InMux I__938 (
            .O(N__5161),
            .I(N__5154));
    InMux I__937 (
            .O(N__5160),
            .I(N__5154));
    InMux I__936 (
            .O(N__5159),
            .I(N__5151));
    LocalMux I__935 (
            .O(N__5154),
            .I(N__5146));
    LocalMux I__934 (
            .O(N__5151),
            .I(N__5146));
    Odrv4 I__933 (
            .O(N__5146),
            .I(r_count_1hzZ0Z_15));
    CascadeMux I__932 (
            .O(N__5143),
            .I(N__5140));
    InMux I__931 (
            .O(N__5140),
            .I(N__5137));
    LocalMux I__930 (
            .O(N__5137),
            .I(N__5134));
    Span4Mux_h I__929 (
            .O(N__5134),
            .I(N__5131));
    Odrv4 I__928 (
            .O(N__5131),
            .I(o_LED_43_4_and));
    InMux I__927 (
            .O(N__5128),
            .I(N__5124));
    InMux I__926 (
            .O(N__5127),
            .I(N__5121));
    LocalMux I__925 (
            .O(N__5124),
            .I(N__5117));
    LocalMux I__924 (
            .O(N__5121),
            .I(N__5113));
    InMux I__923 (
            .O(N__5120),
            .I(N__5110));
    Span4Mux_v I__922 (
            .O(N__5117),
            .I(N__5107));
    InMux I__921 (
            .O(N__5116),
            .I(N__5104));
    Span4Mux_s3_h I__920 (
            .O(N__5113),
            .I(N__5101));
    LocalMux I__919 (
            .O(N__5110),
            .I(r_count_1hzZ0Z_0));
    Odrv4 I__918 (
            .O(N__5107),
            .I(r_count_1hzZ0Z_0));
    LocalMux I__917 (
            .O(N__5104),
            .I(r_count_1hzZ0Z_0));
    Odrv4 I__916 (
            .O(N__5101),
            .I(r_count_1hzZ0Z_0));
    InMux I__915 (
            .O(N__5092),
            .I(N__5089));
    LocalMux I__914 (
            .O(N__5089),
            .I(N__5084));
    CascadeMux I__913 (
            .O(N__5088),
            .I(N__5081));
    InMux I__912 (
            .O(N__5087),
            .I(N__5078));
    Span4Mux_h I__911 (
            .O(N__5084),
            .I(N__5075));
    InMux I__910 (
            .O(N__5081),
            .I(N__5072));
    LocalMux I__909 (
            .O(N__5078),
            .I(r_count_1hzZ0Z_1));
    Odrv4 I__908 (
            .O(N__5075),
            .I(r_count_1hzZ0Z_1));
    LocalMux I__907 (
            .O(N__5072),
            .I(r_count_1hzZ0Z_1));
    CascadeMux I__906 (
            .O(N__5065),
            .I(N__5062));
    InMux I__905 (
            .O(N__5062),
            .I(N__5059));
    LocalMux I__904 (
            .O(N__5059),
            .I(N__5056));
    Span4Mux_h I__903 (
            .O(N__5056),
            .I(N__5052));
    InMux I__902 (
            .O(N__5055),
            .I(N__5049));
    Odrv4 I__901 (
            .O(N__5052),
            .I(r_count_1hzZ0Z_2));
    LocalMux I__900 (
            .O(N__5049),
            .I(r_count_1hzZ0Z_2));
    InMux I__899 (
            .O(N__5044),
            .I(un2_r_count_1hz_1_cry_1));
    InMux I__898 (
            .O(N__5041),
            .I(N__5038));
    LocalMux I__897 (
            .O(N__5038),
            .I(N__5034));
    InMux I__896 (
            .O(N__5037),
            .I(N__5031));
    Span4Mux_h I__895 (
            .O(N__5034),
            .I(N__5028));
    LocalMux I__894 (
            .O(N__5031),
            .I(r_count_1hzZ0Z_3));
    Odrv4 I__893 (
            .O(N__5028),
            .I(r_count_1hzZ0Z_3));
    InMux I__892 (
            .O(N__5023),
            .I(un2_r_count_1hz_1_cry_2));
    InMux I__891 (
            .O(N__5020),
            .I(N__5016));
    InMux I__890 (
            .O(N__5019),
            .I(N__5013));
    LocalMux I__889 (
            .O(N__5016),
            .I(r_count_1hzZ0Z_4));
    LocalMux I__888 (
            .O(N__5013),
            .I(r_count_1hzZ0Z_4));
    InMux I__887 (
            .O(N__5008),
            .I(un2_r_count_1hz_1_cry_3));
    InMux I__886 (
            .O(N__5005),
            .I(N__5002));
    LocalMux I__885 (
            .O(N__5002),
            .I(N__4997));
    InMux I__884 (
            .O(N__5001),
            .I(N__4992));
    InMux I__883 (
            .O(N__5000),
            .I(N__4992));
    Span4Mux_v I__882 (
            .O(N__4997),
            .I(N__4989));
    LocalMux I__881 (
            .O(N__4992),
            .I(r_count_1hzZ0Z_5));
    Odrv4 I__880 (
            .O(N__4989),
            .I(r_count_1hzZ0Z_5));
    InMux I__879 (
            .O(N__4984),
            .I(N__4981));
    LocalMux I__878 (
            .O(N__4981),
            .I(N__4978));
    Span4Mux_v I__877 (
            .O(N__4978),
            .I(N__4975));
    Odrv4 I__876 (
            .O(N__4975),
            .I(un2_r_count_1hz_1_cry_4_THRU_CO));
    InMux I__875 (
            .O(N__4972),
            .I(un2_r_count_1hz_1_cry_4));
    InMux I__874 (
            .O(N__4969),
            .I(N__4965));
    InMux I__873 (
            .O(N__4968),
            .I(N__4962));
    LocalMux I__872 (
            .O(N__4965),
            .I(r_count_1hzZ0Z_6));
    LocalMux I__871 (
            .O(N__4962),
            .I(r_count_1hzZ0Z_6));
    InMux I__870 (
            .O(N__4957),
            .I(un2_r_count_1hz_1_cry_5));
    IoInMux I__869 (
            .O(N__4954),
            .I(N__4951));
    LocalMux I__868 (
            .O(N__4951),
            .I(N__4948));
    Span4Mux_s1_h I__867 (
            .O(N__4948),
            .I(N__4944));
    InMux I__866 (
            .O(N__4947),
            .I(N__4941));
    Odrv4 I__865 (
            .O(N__4944),
            .I(o_LED_1_c));
    LocalMux I__864 (
            .O(N__4941),
            .I(o_LED_1_c));
    CascadeMux I__863 (
            .O(N__4936),
            .I(N__4933));
    InMux I__862 (
            .O(N__4933),
            .I(N__4930));
    LocalMux I__861 (
            .O(N__4930),
            .I(N__4927));
    Odrv12 I__860 (
            .O(N__4927),
            .I(o_LED_13_4_and));
    InMux I__859 (
            .O(N__4924),
            .I(N__4921));
    LocalMux I__858 (
            .O(N__4921),
            .I(N__4918));
    Odrv12 I__857 (
            .O(N__4918),
            .I(o_LED_13_5_and));
    CascadeMux I__856 (
            .O(N__4915),
            .I(N__4912));
    InMux I__855 (
            .O(N__4912),
            .I(N__4909));
    LocalMux I__854 (
            .O(N__4909),
            .I(N__4906));
    Odrv12 I__853 (
            .O(N__4906),
            .I(o_LED_13_6_and));
    CascadeMux I__852 (
            .O(N__4903),
            .I(N__4900));
    InMux I__851 (
            .O(N__4900),
            .I(N__4897));
    LocalMux I__850 (
            .O(N__4897),
            .I(N__4894));
    Odrv12 I__849 (
            .O(N__4894),
            .I(o_LED_13_7_and));
    InMux I__848 (
            .O(N__4891),
            .I(bfn_11_2_0_));
    CascadeMux I__847 (
            .O(N__4888),
            .I(o_LED_13_THRU_CO_cascade_));
    CascadeMux I__846 (
            .O(N__4885),
            .I(N__4882));
    InMux I__845 (
            .O(N__4882),
            .I(N__4879));
    LocalMux I__844 (
            .O(N__4879),
            .I(o_LED_13_1_and));
    CascadeMux I__843 (
            .O(N__4876),
            .I(N__4869));
    CascadeMux I__842 (
            .O(N__4875),
            .I(N__4864));
    CascadeMux I__841 (
            .O(N__4874),
            .I(N__4860));
    CascadeMux I__840 (
            .O(N__4873),
            .I(N__4855));
    InMux I__839 (
            .O(N__4872),
            .I(N__4849));
    InMux I__838 (
            .O(N__4869),
            .I(N__4844));
    InMux I__837 (
            .O(N__4868),
            .I(N__4844));
    InMux I__836 (
            .O(N__4867),
            .I(N__4831));
    InMux I__835 (
            .O(N__4864),
            .I(N__4831));
    InMux I__834 (
            .O(N__4863),
            .I(N__4831));
    InMux I__833 (
            .O(N__4860),
            .I(N__4831));
    InMux I__832 (
            .O(N__4859),
            .I(N__4831));
    InMux I__831 (
            .O(N__4858),
            .I(N__4831));
    InMux I__830 (
            .O(N__4855),
            .I(N__4822));
    InMux I__829 (
            .O(N__4854),
            .I(N__4822));
    InMux I__828 (
            .O(N__4853),
            .I(N__4822));
    InMux I__827 (
            .O(N__4852),
            .I(N__4822));
    LocalMux I__826 (
            .O(N__4849),
            .I(o_LED_43_THRU_CO));
    LocalMux I__825 (
            .O(N__4844),
            .I(o_LED_43_THRU_CO));
    LocalMux I__824 (
            .O(N__4831),
            .I(o_LED_43_THRU_CO));
    LocalMux I__823 (
            .O(N__4822),
            .I(o_LED_43_THRU_CO));
    InMux I__822 (
            .O(N__4813),
            .I(bfn_9_10_0_));
    CascadeMux I__821 (
            .O(N__4810),
            .I(o_LED_43_THRU_CO_cascade_));
    CascadeMux I__820 (
            .O(N__4807),
            .I(N__4804));
    InMux I__819 (
            .O(N__4804),
            .I(N__4801));
    LocalMux I__818 (
            .O(N__4801),
            .I(o_LED_43_1_and));
    CascadeMux I__817 (
            .O(N__4798),
            .I(N__4795));
    InMux I__816 (
            .O(N__4795),
            .I(N__4792));
    LocalMux I__815 (
            .O(N__4792),
            .I(o_LED_43_2_and));
    CascadeMux I__814 (
            .O(N__4789),
            .I(N__4786));
    InMux I__813 (
            .O(N__4786),
            .I(N__4782));
    InMux I__812 (
            .O(N__4785),
            .I(N__4779));
    LocalMux I__811 (
            .O(N__4782),
            .I(N__4776));
    LocalMux I__810 (
            .O(N__4779),
            .I(r_count_5hzZ0Z_28));
    Odrv4 I__809 (
            .O(N__4776),
            .I(r_count_5hzZ0Z_28));
    InMux I__808 (
            .O(N__4771),
            .I(un2_r_count_5hz_1_cry_27));
    InMux I__807 (
            .O(N__4768),
            .I(N__4764));
    InMux I__806 (
            .O(N__4767),
            .I(N__4761));
    LocalMux I__805 (
            .O(N__4764),
            .I(r_count_5hzZ0Z_29));
    LocalMux I__804 (
            .O(N__4761),
            .I(r_count_5hzZ0Z_29));
    InMux I__803 (
            .O(N__4756),
            .I(un2_r_count_5hz_1_cry_28));
    InMux I__802 (
            .O(N__4753),
            .I(N__4749));
    InMux I__801 (
            .O(N__4752),
            .I(N__4746));
    LocalMux I__800 (
            .O(N__4749),
            .I(r_count_5hzZ0Z_30));
    LocalMux I__799 (
            .O(N__4746),
            .I(r_count_5hzZ0Z_30));
    InMux I__798 (
            .O(N__4741),
            .I(un2_r_count_5hz_1_cry_29));
    InMux I__797 (
            .O(N__4738),
            .I(un2_r_count_5hz_1_cry_30));
    InMux I__796 (
            .O(N__4735),
            .I(N__4731));
    InMux I__795 (
            .O(N__4734),
            .I(N__4728));
    LocalMux I__794 (
            .O(N__4731),
            .I(r_count_5hzZ0Z_31));
    LocalMux I__793 (
            .O(N__4728),
            .I(r_count_5hzZ0Z_31));
    CascadeMux I__792 (
            .O(N__4723),
            .I(N__4720));
    InMux I__791 (
            .O(N__4720),
            .I(N__4717));
    LocalMux I__790 (
            .O(N__4717),
            .I(o_LED_43_0_and));
    CascadeMux I__789 (
            .O(N__4714),
            .I(N__4711));
    InMux I__788 (
            .O(N__4711),
            .I(N__4708));
    LocalMux I__787 (
            .O(N__4708),
            .I(o_LED_43_3_and));
    InMux I__786 (
            .O(N__4705),
            .I(N__4701));
    InMux I__785 (
            .O(N__4704),
            .I(N__4698));
    LocalMux I__784 (
            .O(N__4701),
            .I(r_count_5hzZ0Z_20));
    LocalMux I__783 (
            .O(N__4698),
            .I(r_count_5hzZ0Z_20));
    InMux I__782 (
            .O(N__4693),
            .I(un2_r_count_5hz_1_cry_19));
    InMux I__781 (
            .O(N__4690),
            .I(N__4686));
    InMux I__780 (
            .O(N__4689),
            .I(N__4683));
    LocalMux I__779 (
            .O(N__4686),
            .I(N__4680));
    LocalMux I__778 (
            .O(N__4683),
            .I(r_count_5hzZ0Z_21));
    Odrv4 I__777 (
            .O(N__4680),
            .I(r_count_5hzZ0Z_21));
    InMux I__776 (
            .O(N__4675),
            .I(un2_r_count_5hz_1_cry_20));
    CascadeMux I__775 (
            .O(N__4672),
            .I(N__4668));
    InMux I__774 (
            .O(N__4671),
            .I(N__4665));
    InMux I__773 (
            .O(N__4668),
            .I(N__4662));
    LocalMux I__772 (
            .O(N__4665),
            .I(r_count_5hzZ0Z_22));
    LocalMux I__771 (
            .O(N__4662),
            .I(r_count_5hzZ0Z_22));
    InMux I__770 (
            .O(N__4657),
            .I(un2_r_count_5hz_1_cry_21));
    InMux I__769 (
            .O(N__4654),
            .I(N__4650));
    InMux I__768 (
            .O(N__4653),
            .I(N__4647));
    LocalMux I__767 (
            .O(N__4650),
            .I(N__4642));
    LocalMux I__766 (
            .O(N__4647),
            .I(N__4642));
    Odrv4 I__765 (
            .O(N__4642),
            .I(r_count_5hzZ0Z_23));
    InMux I__764 (
            .O(N__4639),
            .I(un2_r_count_5hz_1_cry_22));
    InMux I__763 (
            .O(N__4636),
            .I(N__4632));
    InMux I__762 (
            .O(N__4635),
            .I(N__4629));
    LocalMux I__761 (
            .O(N__4632),
            .I(r_count_5hzZ0Z_24));
    LocalMux I__760 (
            .O(N__4629),
            .I(r_count_5hzZ0Z_24));
    InMux I__759 (
            .O(N__4624),
            .I(un2_r_count_5hz_1_cry_23));
    InMux I__758 (
            .O(N__4621),
            .I(N__4617));
    InMux I__757 (
            .O(N__4620),
            .I(N__4614));
    LocalMux I__756 (
            .O(N__4617),
            .I(r_count_5hzZ0Z_25));
    LocalMux I__755 (
            .O(N__4614),
            .I(r_count_5hzZ0Z_25));
    InMux I__754 (
            .O(N__4609),
            .I(bfn_9_5_0_));
    CascadeMux I__753 (
            .O(N__4606),
            .I(N__4602));
    InMux I__752 (
            .O(N__4605),
            .I(N__4599));
    InMux I__751 (
            .O(N__4602),
            .I(N__4596));
    LocalMux I__750 (
            .O(N__4599),
            .I(r_count_5hzZ0Z_26));
    LocalMux I__749 (
            .O(N__4596),
            .I(r_count_5hzZ0Z_26));
    InMux I__748 (
            .O(N__4591),
            .I(un2_r_count_5hz_1_cry_25));
    InMux I__747 (
            .O(N__4588),
            .I(N__4584));
    InMux I__746 (
            .O(N__4587),
            .I(N__4581));
    LocalMux I__745 (
            .O(N__4584),
            .I(r_count_5hzZ0Z_27));
    LocalMux I__744 (
            .O(N__4581),
            .I(r_count_5hzZ0Z_27));
    InMux I__743 (
            .O(N__4576),
            .I(un2_r_count_5hz_1_cry_26));
    InMux I__742 (
            .O(N__4573),
            .I(N__4568));
    InMux I__741 (
            .O(N__4572),
            .I(N__4563));
    InMux I__740 (
            .O(N__4571),
            .I(N__4563));
    LocalMux I__739 (
            .O(N__4568),
            .I(r_count_5hzZ0Z_12));
    LocalMux I__738 (
            .O(N__4563),
            .I(r_count_5hzZ0Z_12));
    InMux I__737 (
            .O(N__4558),
            .I(N__4555));
    LocalMux I__736 (
            .O(N__4555),
            .I(un2_r_count_5hz_1_cry_11_THRU_CO));
    InMux I__735 (
            .O(N__4552),
            .I(un2_r_count_5hz_1_cry_11));
    InMux I__734 (
            .O(N__4549),
            .I(N__4545));
    InMux I__733 (
            .O(N__4548),
            .I(N__4542));
    LocalMux I__732 (
            .O(N__4545),
            .I(r_count_5hzZ0Z_13));
    LocalMux I__731 (
            .O(N__4542),
            .I(r_count_5hzZ0Z_13));
    InMux I__730 (
            .O(N__4537),
            .I(un2_r_count_5hz_1_cry_12));
    CascadeMux I__729 (
            .O(N__4534),
            .I(N__4529));
    InMux I__728 (
            .O(N__4533),
            .I(N__4526));
    InMux I__727 (
            .O(N__4532),
            .I(N__4523));
    InMux I__726 (
            .O(N__4529),
            .I(N__4520));
    LocalMux I__725 (
            .O(N__4526),
            .I(r_count_5hzZ0Z_14));
    LocalMux I__724 (
            .O(N__4523),
            .I(r_count_5hzZ0Z_14));
    LocalMux I__723 (
            .O(N__4520),
            .I(r_count_5hzZ0Z_14));
    InMux I__722 (
            .O(N__4513),
            .I(N__4510));
    LocalMux I__721 (
            .O(N__4510),
            .I(un2_r_count_5hz_1_cry_13_THRU_CO));
    InMux I__720 (
            .O(N__4507),
            .I(un2_r_count_5hz_1_cry_13));
    InMux I__719 (
            .O(N__4504),
            .I(N__4499));
    InMux I__718 (
            .O(N__4503),
            .I(N__4494));
    InMux I__717 (
            .O(N__4502),
            .I(N__4494));
    LocalMux I__716 (
            .O(N__4499),
            .I(r_count_5hzZ0Z_15));
    LocalMux I__715 (
            .O(N__4494),
            .I(r_count_5hzZ0Z_15));
    InMux I__714 (
            .O(N__4489),
            .I(N__4486));
    LocalMux I__713 (
            .O(N__4486),
            .I(un2_r_count_5hz_1_cry_14_THRU_CO));
    InMux I__712 (
            .O(N__4483),
            .I(un2_r_count_5hz_1_cry_14));
    InMux I__711 (
            .O(N__4480),
            .I(N__4475));
    InMux I__710 (
            .O(N__4479),
            .I(N__4472));
    InMux I__709 (
            .O(N__4478),
            .I(N__4469));
    LocalMux I__708 (
            .O(N__4475),
            .I(N__4466));
    LocalMux I__707 (
            .O(N__4472),
            .I(r_count_5hzZ0Z_16));
    LocalMux I__706 (
            .O(N__4469),
            .I(r_count_5hzZ0Z_16));
    Odrv4 I__705 (
            .O(N__4466),
            .I(r_count_5hzZ0Z_16));
    InMux I__704 (
            .O(N__4459),
            .I(N__4456));
    LocalMux I__703 (
            .O(N__4456),
            .I(un2_r_count_5hz_1_cry_15_THRU_CO));
    InMux I__702 (
            .O(N__4453),
            .I(un2_r_count_5hz_1_cry_15));
    InMux I__701 (
            .O(N__4450),
            .I(N__4445));
    InMux I__700 (
            .O(N__4449),
            .I(N__4442));
    InMux I__699 (
            .O(N__4448),
            .I(N__4439));
    LocalMux I__698 (
            .O(N__4445),
            .I(r_count_5hzZ0Z_17));
    LocalMux I__697 (
            .O(N__4442),
            .I(r_count_5hzZ0Z_17));
    LocalMux I__696 (
            .O(N__4439),
            .I(r_count_5hzZ0Z_17));
    InMux I__695 (
            .O(N__4432),
            .I(N__4429));
    LocalMux I__694 (
            .O(N__4429),
            .I(un2_r_count_5hz_1_cry_16_THRU_CO));
    InMux I__693 (
            .O(N__4426),
            .I(bfn_9_4_0_));
    CascadeMux I__692 (
            .O(N__4423),
            .I(N__4419));
    InMux I__691 (
            .O(N__4422),
            .I(N__4416));
    InMux I__690 (
            .O(N__4419),
            .I(N__4413));
    LocalMux I__689 (
            .O(N__4416),
            .I(N__4408));
    LocalMux I__688 (
            .O(N__4413),
            .I(N__4408));
    Odrv4 I__687 (
            .O(N__4408),
            .I(r_count_5hzZ0Z_18));
    InMux I__686 (
            .O(N__4405),
            .I(un2_r_count_5hz_1_cry_17));
    InMux I__685 (
            .O(N__4402),
            .I(N__4398));
    InMux I__684 (
            .O(N__4401),
            .I(N__4395));
    LocalMux I__683 (
            .O(N__4398),
            .I(r_count_5hzZ0Z_19));
    LocalMux I__682 (
            .O(N__4395),
            .I(r_count_5hzZ0Z_19));
    InMux I__681 (
            .O(N__4390),
            .I(un2_r_count_5hz_1_cry_18));
    InMux I__680 (
            .O(N__4387),
            .I(N__4380));
    InMux I__679 (
            .O(N__4386),
            .I(N__4380));
    InMux I__678 (
            .O(N__4385),
            .I(N__4377));
    LocalMux I__677 (
            .O(N__4380),
            .I(r_count_5hzZ0Z_4));
    LocalMux I__676 (
            .O(N__4377),
            .I(r_count_5hzZ0Z_4));
    InMux I__675 (
            .O(N__4372),
            .I(N__4369));
    LocalMux I__674 (
            .O(N__4369),
            .I(un2_r_count_5hz_1_cry_3_THRU_CO));
    InMux I__673 (
            .O(N__4366),
            .I(un2_r_count_5hz_1_cry_3));
    InMux I__672 (
            .O(N__4363),
            .I(N__4359));
    InMux I__671 (
            .O(N__4362),
            .I(N__4356));
    LocalMux I__670 (
            .O(N__4359),
            .I(r_count_5hzZ0Z_5));
    LocalMux I__669 (
            .O(N__4356),
            .I(r_count_5hzZ0Z_5));
    InMux I__668 (
            .O(N__4351),
            .I(un2_r_count_5hz_1_cry_4));
    CascadeMux I__667 (
            .O(N__4348),
            .I(N__4345));
    InMux I__666 (
            .O(N__4345),
            .I(N__4341));
    InMux I__665 (
            .O(N__4344),
            .I(N__4338));
    LocalMux I__664 (
            .O(N__4341),
            .I(r_count_5hzZ0Z_6));
    LocalMux I__663 (
            .O(N__4338),
            .I(r_count_5hzZ0Z_6));
    InMux I__662 (
            .O(N__4333),
            .I(un2_r_count_5hz_1_cry_5));
    InMux I__661 (
            .O(N__4330),
            .I(N__4325));
    InMux I__660 (
            .O(N__4329),
            .I(N__4322));
    InMux I__659 (
            .O(N__4328),
            .I(N__4319));
    LocalMux I__658 (
            .O(N__4325),
            .I(r_count_5hzZ0Z_7));
    LocalMux I__657 (
            .O(N__4322),
            .I(r_count_5hzZ0Z_7));
    LocalMux I__656 (
            .O(N__4319),
            .I(r_count_5hzZ0Z_7));
    InMux I__655 (
            .O(N__4312),
            .I(N__4309));
    LocalMux I__654 (
            .O(N__4309),
            .I(un2_r_count_5hz_1_cry_6_THRU_CO));
    InMux I__653 (
            .O(N__4306),
            .I(un2_r_count_5hz_1_cry_6));
    InMux I__652 (
            .O(N__4303),
            .I(N__4299));
    InMux I__651 (
            .O(N__4302),
            .I(N__4296));
    LocalMux I__650 (
            .O(N__4299),
            .I(r_count_5hzZ0Z_8));
    LocalMux I__649 (
            .O(N__4296),
            .I(r_count_5hzZ0Z_8));
    InMux I__648 (
            .O(N__4291),
            .I(un2_r_count_5hz_1_cry_7));
    InMux I__647 (
            .O(N__4288),
            .I(N__4284));
    InMux I__646 (
            .O(N__4287),
            .I(N__4281));
    LocalMux I__645 (
            .O(N__4284),
            .I(r_count_5hzZ0Z_9));
    LocalMux I__644 (
            .O(N__4281),
            .I(r_count_5hzZ0Z_9));
    InMux I__643 (
            .O(N__4276),
            .I(bfn_9_3_0_));
    InMux I__642 (
            .O(N__4273),
            .I(N__4269));
    InMux I__641 (
            .O(N__4272),
            .I(N__4266));
    LocalMux I__640 (
            .O(N__4269),
            .I(r_count_5hzZ0Z_10));
    LocalMux I__639 (
            .O(N__4266),
            .I(r_count_5hzZ0Z_10));
    InMux I__638 (
            .O(N__4261),
            .I(un2_r_count_5hz_1_cry_9));
    InMux I__637 (
            .O(N__4258),
            .I(N__4254));
    InMux I__636 (
            .O(N__4257),
            .I(N__4251));
    LocalMux I__635 (
            .O(N__4254),
            .I(r_count_5hzZ0Z_11));
    LocalMux I__634 (
            .O(N__4251),
            .I(r_count_5hzZ0Z_11));
    InMux I__633 (
            .O(N__4246),
            .I(un2_r_count_5hz_1_cry_10));
    InMux I__632 (
            .O(N__4243),
            .I(un2_r_count_2hz_1_cry_30));
    InMux I__631 (
            .O(N__4240),
            .I(N__4236));
    InMux I__630 (
            .O(N__4239),
            .I(N__4233));
    LocalMux I__629 (
            .O(N__4236),
            .I(r_count_2hzZ0Z_31));
    LocalMux I__628 (
            .O(N__4233),
            .I(r_count_2hzZ0Z_31));
    IoInMux I__627 (
            .O(N__4228),
            .I(N__4225));
    LocalMux I__626 (
            .O(N__4225),
            .I(N__4222));
    Span4Mux_s3_h I__625 (
            .O(N__4222),
            .I(N__4218));
    InMux I__624 (
            .O(N__4221),
            .I(N__4215));
    Odrv4 I__623 (
            .O(N__4218),
            .I(o_LED_4_c));
    LocalMux I__622 (
            .O(N__4215),
            .I(o_LED_4_c));
    CascadeMux I__621 (
            .O(N__4210),
            .I(N__4205));
    InMux I__620 (
            .O(N__4209),
            .I(N__4201));
    InMux I__619 (
            .O(N__4208),
            .I(N__4196));
    InMux I__618 (
            .O(N__4205),
            .I(N__4196));
    InMux I__617 (
            .O(N__4204),
            .I(N__4193));
    LocalMux I__616 (
            .O(N__4201),
            .I(r_count_5hzZ0Z_0));
    LocalMux I__615 (
            .O(N__4196),
            .I(r_count_5hzZ0Z_0));
    LocalMux I__614 (
            .O(N__4193),
            .I(r_count_5hzZ0Z_0));
    CascadeMux I__613 (
            .O(N__4186),
            .I(N__4181));
    InMux I__612 (
            .O(N__4185),
            .I(N__4176));
    InMux I__611 (
            .O(N__4184),
            .I(N__4176));
    InMux I__610 (
            .O(N__4181),
            .I(N__4173));
    LocalMux I__609 (
            .O(N__4176),
            .I(r_count_5hzZ0Z_1));
    LocalMux I__608 (
            .O(N__4173),
            .I(r_count_5hzZ0Z_1));
    InMux I__607 (
            .O(N__4168),
            .I(N__4165));
    LocalMux I__606 (
            .O(N__4165),
            .I(N__4161));
    InMux I__605 (
            .O(N__4164),
            .I(N__4158));
    Odrv4 I__604 (
            .O(N__4161),
            .I(r_count_5hzZ0Z_2));
    LocalMux I__603 (
            .O(N__4158),
            .I(r_count_5hzZ0Z_2));
    InMux I__602 (
            .O(N__4153),
            .I(un2_r_count_5hz_1_cry_1));
    CascadeMux I__601 (
            .O(N__4150),
            .I(N__4147));
    InMux I__600 (
            .O(N__4147),
            .I(N__4143));
    InMux I__599 (
            .O(N__4146),
            .I(N__4140));
    LocalMux I__598 (
            .O(N__4143),
            .I(r_count_5hzZ0Z_3));
    LocalMux I__597 (
            .O(N__4140),
            .I(r_count_5hzZ0Z_3));
    InMux I__596 (
            .O(N__4135),
            .I(un2_r_count_5hz_1_cry_2));
    CascadeMux I__595 (
            .O(N__4132),
            .I(N__4127));
    InMux I__594 (
            .O(N__4131),
            .I(N__4124));
    InMux I__593 (
            .O(N__4130),
            .I(N__4121));
    InMux I__592 (
            .O(N__4127),
            .I(N__4118));
    LocalMux I__591 (
            .O(N__4124),
            .I(r_count_2hzZ0Z_22));
    LocalMux I__590 (
            .O(N__4121),
            .I(r_count_2hzZ0Z_22));
    LocalMux I__589 (
            .O(N__4118),
            .I(r_count_2hzZ0Z_22));
    InMux I__588 (
            .O(N__4111),
            .I(N__4108));
    LocalMux I__587 (
            .O(N__4108),
            .I(un2_r_count_2hz_1_cry_21_THRU_CO));
    InMux I__586 (
            .O(N__4105),
            .I(un2_r_count_2hz_1_cry_21));
    InMux I__585 (
            .O(N__4102),
            .I(N__4098));
    InMux I__584 (
            .O(N__4101),
            .I(N__4095));
    LocalMux I__583 (
            .O(N__4098),
            .I(r_count_2hzZ0Z_23));
    LocalMux I__582 (
            .O(N__4095),
            .I(r_count_2hzZ0Z_23));
    InMux I__581 (
            .O(N__4090),
            .I(un2_r_count_2hz_1_cry_22));
    CascadeMux I__580 (
            .O(N__4087),
            .I(N__4083));
    InMux I__579 (
            .O(N__4086),
            .I(N__4080));
    InMux I__578 (
            .O(N__4083),
            .I(N__4077));
    LocalMux I__577 (
            .O(N__4080),
            .I(r_count_2hzZ0Z_24));
    LocalMux I__576 (
            .O(N__4077),
            .I(r_count_2hzZ0Z_24));
    InMux I__575 (
            .O(N__4072),
            .I(un2_r_count_2hz_1_cry_23));
    InMux I__574 (
            .O(N__4069),
            .I(N__4065));
    InMux I__573 (
            .O(N__4068),
            .I(N__4062));
    LocalMux I__572 (
            .O(N__4065),
            .I(r_count_2hzZ0Z_25));
    LocalMux I__571 (
            .O(N__4062),
            .I(r_count_2hzZ0Z_25));
    InMux I__570 (
            .O(N__4057),
            .I(bfn_8_9_0_));
    InMux I__569 (
            .O(N__4054),
            .I(N__4050));
    InMux I__568 (
            .O(N__4053),
            .I(N__4047));
    LocalMux I__567 (
            .O(N__4050),
            .I(N__4044));
    LocalMux I__566 (
            .O(N__4047),
            .I(r_count_2hzZ0Z_26));
    Odrv4 I__565 (
            .O(N__4044),
            .I(r_count_2hzZ0Z_26));
    InMux I__564 (
            .O(N__4039),
            .I(un2_r_count_2hz_1_cry_25));
    InMux I__563 (
            .O(N__4036),
            .I(N__4032));
    InMux I__562 (
            .O(N__4035),
            .I(N__4029));
    LocalMux I__561 (
            .O(N__4032),
            .I(r_count_2hzZ0Z_27));
    LocalMux I__560 (
            .O(N__4029),
            .I(r_count_2hzZ0Z_27));
    InMux I__559 (
            .O(N__4024),
            .I(un2_r_count_2hz_1_cry_26));
    InMux I__558 (
            .O(N__4021),
            .I(N__4017));
    InMux I__557 (
            .O(N__4020),
            .I(N__4014));
    LocalMux I__556 (
            .O(N__4017),
            .I(r_count_2hzZ0Z_28));
    LocalMux I__555 (
            .O(N__4014),
            .I(r_count_2hzZ0Z_28));
    InMux I__554 (
            .O(N__4009),
            .I(un2_r_count_2hz_1_cry_27));
    InMux I__553 (
            .O(N__4006),
            .I(N__4002));
    InMux I__552 (
            .O(N__4005),
            .I(N__3999));
    LocalMux I__551 (
            .O(N__4002),
            .I(r_count_2hzZ0Z_29));
    LocalMux I__550 (
            .O(N__3999),
            .I(r_count_2hzZ0Z_29));
    InMux I__549 (
            .O(N__3994),
            .I(un2_r_count_2hz_1_cry_28));
    CascadeMux I__548 (
            .O(N__3991),
            .I(N__3987));
    InMux I__547 (
            .O(N__3990),
            .I(N__3984));
    InMux I__546 (
            .O(N__3987),
            .I(N__3981));
    LocalMux I__545 (
            .O(N__3984),
            .I(r_count_2hzZ0Z_30));
    LocalMux I__544 (
            .O(N__3981),
            .I(r_count_2hzZ0Z_30));
    InMux I__543 (
            .O(N__3976),
            .I(un2_r_count_2hz_1_cry_29));
    InMux I__542 (
            .O(N__3973),
            .I(N__3970));
    LocalMux I__541 (
            .O(N__3970),
            .I(N__3965));
    InMux I__540 (
            .O(N__3969),
            .I(N__3962));
    InMux I__539 (
            .O(N__3968),
            .I(N__3959));
    Odrv4 I__538 (
            .O(N__3965),
            .I(r_count_2hzZ0Z_14));
    LocalMux I__537 (
            .O(N__3962),
            .I(r_count_2hzZ0Z_14));
    LocalMux I__536 (
            .O(N__3959),
            .I(r_count_2hzZ0Z_14));
    InMux I__535 (
            .O(N__3952),
            .I(N__3949));
    LocalMux I__534 (
            .O(N__3949),
            .I(un2_r_count_2hz_1_cry_13_THRU_CO));
    InMux I__533 (
            .O(N__3946),
            .I(un2_r_count_2hz_1_cry_13));
    CascadeMux I__532 (
            .O(N__3943),
            .I(N__3939));
    InMux I__531 (
            .O(N__3942),
            .I(N__3936));
    InMux I__530 (
            .O(N__3939),
            .I(N__3933));
    LocalMux I__529 (
            .O(N__3936),
            .I(r_count_2hzZ0Z_15));
    LocalMux I__528 (
            .O(N__3933),
            .I(r_count_2hzZ0Z_15));
    InMux I__527 (
            .O(N__3928),
            .I(un2_r_count_2hz_1_cry_14));
    InMux I__526 (
            .O(N__3925),
            .I(N__3920));
    InMux I__525 (
            .O(N__3924),
            .I(N__3917));
    InMux I__524 (
            .O(N__3923),
            .I(N__3914));
    LocalMux I__523 (
            .O(N__3920),
            .I(r_count_2hzZ0Z_16));
    LocalMux I__522 (
            .O(N__3917),
            .I(r_count_2hzZ0Z_16));
    LocalMux I__521 (
            .O(N__3914),
            .I(r_count_2hzZ0Z_16));
    InMux I__520 (
            .O(N__3907),
            .I(N__3904));
    LocalMux I__519 (
            .O(N__3904),
            .I(N__3901));
    Odrv4 I__518 (
            .O(N__3901),
            .I(un2_r_count_2hz_1_cry_15_THRU_CO));
    InMux I__517 (
            .O(N__3898),
            .I(un2_r_count_2hz_1_cry_15));
    InMux I__516 (
            .O(N__3895),
            .I(N__3892));
    LocalMux I__515 (
            .O(N__3892),
            .I(N__3887));
    InMux I__514 (
            .O(N__3891),
            .I(N__3882));
    InMux I__513 (
            .O(N__3890),
            .I(N__3882));
    Odrv4 I__512 (
            .O(N__3887),
            .I(r_count_2hzZ0Z_17));
    LocalMux I__511 (
            .O(N__3882),
            .I(r_count_2hzZ0Z_17));
    InMux I__510 (
            .O(N__3877),
            .I(N__3874));
    LocalMux I__509 (
            .O(N__3874),
            .I(N__3871));
    Odrv4 I__508 (
            .O(N__3871),
            .I(un2_r_count_2hz_1_cry_16_THRU_CO));
    InMux I__507 (
            .O(N__3868),
            .I(bfn_8_8_0_));
    InMux I__506 (
            .O(N__3865),
            .I(N__3860));
    InMux I__505 (
            .O(N__3864),
            .I(N__3857));
    InMux I__504 (
            .O(N__3863),
            .I(N__3854));
    LocalMux I__503 (
            .O(N__3860),
            .I(r_count_2hzZ0Z_18));
    LocalMux I__502 (
            .O(N__3857),
            .I(r_count_2hzZ0Z_18));
    LocalMux I__501 (
            .O(N__3854),
            .I(r_count_2hzZ0Z_18));
    InMux I__500 (
            .O(N__3847),
            .I(N__3844));
    LocalMux I__499 (
            .O(N__3844),
            .I(un2_r_count_2hz_1_cry_17_THRU_CO));
    InMux I__498 (
            .O(N__3841),
            .I(un2_r_count_2hz_1_cry_17));
    InMux I__497 (
            .O(N__3838),
            .I(N__3833));
    InMux I__496 (
            .O(N__3837),
            .I(N__3830));
    InMux I__495 (
            .O(N__3836),
            .I(N__3827));
    LocalMux I__494 (
            .O(N__3833),
            .I(r_count_2hzZ0Z_19));
    LocalMux I__493 (
            .O(N__3830),
            .I(r_count_2hzZ0Z_19));
    LocalMux I__492 (
            .O(N__3827),
            .I(r_count_2hzZ0Z_19));
    InMux I__491 (
            .O(N__3820),
            .I(N__3817));
    LocalMux I__490 (
            .O(N__3817),
            .I(N__3814));
    Odrv4 I__489 (
            .O(N__3814),
            .I(un2_r_count_2hz_1_cry_18_THRU_CO));
    InMux I__488 (
            .O(N__3811),
            .I(un2_r_count_2hz_1_cry_18));
    InMux I__487 (
            .O(N__3808),
            .I(N__3803));
    InMux I__486 (
            .O(N__3807),
            .I(N__3800));
    InMux I__485 (
            .O(N__3806),
            .I(N__3797));
    LocalMux I__484 (
            .O(N__3803),
            .I(r_count_2hzZ0Z_20));
    LocalMux I__483 (
            .O(N__3800),
            .I(r_count_2hzZ0Z_20));
    LocalMux I__482 (
            .O(N__3797),
            .I(r_count_2hzZ0Z_20));
    InMux I__481 (
            .O(N__3790),
            .I(N__3787));
    LocalMux I__480 (
            .O(N__3787),
            .I(un2_r_count_2hz_1_cry_19_THRU_CO));
    InMux I__479 (
            .O(N__3784),
            .I(un2_r_count_2hz_1_cry_19));
    InMux I__478 (
            .O(N__3781),
            .I(N__3777));
    InMux I__477 (
            .O(N__3780),
            .I(N__3774));
    LocalMux I__476 (
            .O(N__3777),
            .I(r_count_2hzZ0Z_21));
    LocalMux I__475 (
            .O(N__3774),
            .I(r_count_2hzZ0Z_21));
    InMux I__474 (
            .O(N__3769),
            .I(un2_r_count_2hz_1_cry_20));
    InMux I__473 (
            .O(N__3766),
            .I(N__3762));
    InMux I__472 (
            .O(N__3765),
            .I(N__3759));
    LocalMux I__471 (
            .O(N__3762),
            .I(r_count_2hzZ0Z_6));
    LocalMux I__470 (
            .O(N__3759),
            .I(r_count_2hzZ0Z_6));
    InMux I__469 (
            .O(N__3754),
            .I(un2_r_count_2hz_1_cry_5));
    CascadeMux I__468 (
            .O(N__3751),
            .I(N__3748));
    InMux I__467 (
            .O(N__3748),
            .I(N__3744));
    InMux I__466 (
            .O(N__3747),
            .I(N__3741));
    LocalMux I__465 (
            .O(N__3744),
            .I(r_count_2hzZ0Z_7));
    LocalMux I__464 (
            .O(N__3741),
            .I(r_count_2hzZ0Z_7));
    InMux I__463 (
            .O(N__3736),
            .I(un2_r_count_2hz_1_cry_6));
    InMux I__462 (
            .O(N__3733),
            .I(N__3729));
    InMux I__461 (
            .O(N__3732),
            .I(N__3726));
    LocalMux I__460 (
            .O(N__3729),
            .I(r_count_2hzZ0Z_8));
    LocalMux I__459 (
            .O(N__3726),
            .I(r_count_2hzZ0Z_8));
    InMux I__458 (
            .O(N__3721),
            .I(un2_r_count_2hz_1_cry_7));
    CascadeMux I__457 (
            .O(N__3718),
            .I(N__3715));
    InMux I__456 (
            .O(N__3715),
            .I(N__3708));
    InMux I__455 (
            .O(N__3714),
            .I(N__3708));
    InMux I__454 (
            .O(N__3713),
            .I(N__3705));
    LocalMux I__453 (
            .O(N__3708),
            .I(r_count_2hzZ0Z_9));
    LocalMux I__452 (
            .O(N__3705),
            .I(r_count_2hzZ0Z_9));
    InMux I__451 (
            .O(N__3700),
            .I(N__3697));
    LocalMux I__450 (
            .O(N__3697),
            .I(un2_r_count_2hz_1_cry_8_THRU_CO));
    InMux I__449 (
            .O(N__3694),
            .I(bfn_8_7_0_));
    CascadeMux I__448 (
            .O(N__3691),
            .I(N__3687));
    CascadeMux I__447 (
            .O(N__3690),
            .I(N__3684));
    InMux I__446 (
            .O(N__3687),
            .I(N__3678));
    InMux I__445 (
            .O(N__3684),
            .I(N__3678));
    InMux I__444 (
            .O(N__3683),
            .I(N__3675));
    LocalMux I__443 (
            .O(N__3678),
            .I(N__3672));
    LocalMux I__442 (
            .O(N__3675),
            .I(r_count_2hzZ0Z_10));
    Odrv4 I__441 (
            .O(N__3672),
            .I(r_count_2hzZ0Z_10));
    InMux I__440 (
            .O(N__3667),
            .I(N__3664));
    LocalMux I__439 (
            .O(N__3664),
            .I(un2_r_count_2hz_1_cry_9_THRU_CO));
    InMux I__438 (
            .O(N__3661),
            .I(un2_r_count_2hz_1_cry_9));
    InMux I__437 (
            .O(N__3658),
            .I(N__3653));
    InMux I__436 (
            .O(N__3657),
            .I(N__3648));
    InMux I__435 (
            .O(N__3656),
            .I(N__3648));
    LocalMux I__434 (
            .O(N__3653),
            .I(r_count_2hzZ0Z_11));
    LocalMux I__433 (
            .O(N__3648),
            .I(r_count_2hzZ0Z_11));
    InMux I__432 (
            .O(N__3643),
            .I(N__3640));
    LocalMux I__431 (
            .O(N__3640),
            .I(un2_r_count_2hz_1_cry_10_THRU_CO));
    InMux I__430 (
            .O(N__3637),
            .I(un2_r_count_2hz_1_cry_10));
    CascadeMux I__429 (
            .O(N__3634),
            .I(N__3629));
    InMux I__428 (
            .O(N__3633),
            .I(N__3626));
    InMux I__427 (
            .O(N__3632),
            .I(N__3623));
    InMux I__426 (
            .O(N__3629),
            .I(N__3620));
    LocalMux I__425 (
            .O(N__3626),
            .I(r_count_2hzZ0Z_12));
    LocalMux I__424 (
            .O(N__3623),
            .I(r_count_2hzZ0Z_12));
    LocalMux I__423 (
            .O(N__3620),
            .I(r_count_2hzZ0Z_12));
    InMux I__422 (
            .O(N__3613),
            .I(N__3610));
    LocalMux I__421 (
            .O(N__3610),
            .I(un2_r_count_2hz_1_cry_11_THRU_CO));
    InMux I__420 (
            .O(N__3607),
            .I(un2_r_count_2hz_1_cry_11));
    InMux I__419 (
            .O(N__3604),
            .I(N__3600));
    InMux I__418 (
            .O(N__3603),
            .I(N__3597));
    LocalMux I__417 (
            .O(N__3600),
            .I(r_count_2hzZ0Z_13));
    LocalMux I__416 (
            .O(N__3597),
            .I(r_count_2hzZ0Z_13));
    InMux I__415 (
            .O(N__3592),
            .I(un2_r_count_2hz_1_cry_12));
    CascadeMux I__414 (
            .O(N__3589),
            .I(N__3586));
    InMux I__413 (
            .O(N__3586),
            .I(N__3583));
    LocalMux I__412 (
            .O(N__3583),
            .I(o_LED_23_6_and));
    CascadeMux I__411 (
            .O(N__3580),
            .I(N__3577));
    InMux I__410 (
            .O(N__3577),
            .I(N__3574));
    LocalMux I__409 (
            .O(N__3574),
            .I(o_LED_23_4_and));
    CascadeMux I__408 (
            .O(N__3571),
            .I(N__3564));
    CascadeMux I__407 (
            .O(N__3570),
            .I(N__3560));
    CascadeMux I__406 (
            .O(N__3569),
            .I(N__3555));
    CascadeMux I__405 (
            .O(N__3568),
            .I(N__3551));
    InMux I__404 (
            .O(N__3567),
            .I(N__3538));
    InMux I__403 (
            .O(N__3564),
            .I(N__3538));
    InMux I__402 (
            .O(N__3563),
            .I(N__3538));
    InMux I__401 (
            .O(N__3560),
            .I(N__3538));
    InMux I__400 (
            .O(N__3559),
            .I(N__3538));
    InMux I__399 (
            .O(N__3558),
            .I(N__3538));
    InMux I__398 (
            .O(N__3555),
            .I(N__3531));
    InMux I__397 (
            .O(N__3554),
            .I(N__3531));
    InMux I__396 (
            .O(N__3551),
            .I(N__3531));
    LocalMux I__395 (
            .O(N__3538),
            .I(o_LED_23_THRU_CO));
    LocalMux I__394 (
            .O(N__3531),
            .I(o_LED_23_THRU_CO));
    InMux I__393 (
            .O(N__3526),
            .I(N__3520));
    InMux I__392 (
            .O(N__3525),
            .I(N__3515));
    InMux I__391 (
            .O(N__3524),
            .I(N__3515));
    InMux I__390 (
            .O(N__3523),
            .I(N__3512));
    LocalMux I__389 (
            .O(N__3520),
            .I(r_count_2hzZ0Z_0));
    LocalMux I__388 (
            .O(N__3515),
            .I(r_count_2hzZ0Z_0));
    LocalMux I__387 (
            .O(N__3512),
            .I(r_count_2hzZ0Z_0));
    CascadeMux I__386 (
            .O(N__3505),
            .I(N__3500));
    InMux I__385 (
            .O(N__3504),
            .I(N__3497));
    InMux I__384 (
            .O(N__3503),
            .I(N__3494));
    InMux I__383 (
            .O(N__3500),
            .I(N__3491));
    LocalMux I__382 (
            .O(N__3497),
            .I(r_count_2hzZ0Z_1));
    LocalMux I__381 (
            .O(N__3494),
            .I(r_count_2hzZ0Z_1));
    LocalMux I__380 (
            .O(N__3491),
            .I(r_count_2hzZ0Z_1));
    CascadeMux I__379 (
            .O(N__3484),
            .I(N__3480));
    InMux I__378 (
            .O(N__3483),
            .I(N__3477));
    InMux I__377 (
            .O(N__3480),
            .I(N__3474));
    LocalMux I__376 (
            .O(N__3477),
            .I(r_count_2hzZ0Z_2));
    LocalMux I__375 (
            .O(N__3474),
            .I(r_count_2hzZ0Z_2));
    InMux I__374 (
            .O(N__3469),
            .I(un2_r_count_2hz_1_cry_1));
    InMux I__373 (
            .O(N__3466),
            .I(N__3462));
    InMux I__372 (
            .O(N__3465),
            .I(N__3459));
    LocalMux I__371 (
            .O(N__3462),
            .I(r_count_2hzZ0Z_3));
    LocalMux I__370 (
            .O(N__3459),
            .I(r_count_2hzZ0Z_3));
    InMux I__369 (
            .O(N__3454),
            .I(un2_r_count_2hz_1_cry_2));
    InMux I__368 (
            .O(N__3451),
            .I(N__3444));
    InMux I__367 (
            .O(N__3450),
            .I(N__3444));
    InMux I__366 (
            .O(N__3449),
            .I(N__3441));
    LocalMux I__365 (
            .O(N__3444),
            .I(r_count_2hzZ0Z_4));
    LocalMux I__364 (
            .O(N__3441),
            .I(r_count_2hzZ0Z_4));
    InMux I__363 (
            .O(N__3436),
            .I(N__3433));
    LocalMux I__362 (
            .O(N__3433),
            .I(un2_r_count_2hz_1_cry_3_THRU_CO));
    InMux I__361 (
            .O(N__3430),
            .I(un2_r_count_2hz_1_cry_3));
    InMux I__360 (
            .O(N__3427),
            .I(N__3423));
    InMux I__359 (
            .O(N__3426),
            .I(N__3420));
    LocalMux I__358 (
            .O(N__3423),
            .I(r_count_2hzZ0Z_5));
    LocalMux I__357 (
            .O(N__3420),
            .I(r_count_2hzZ0Z_5));
    InMux I__356 (
            .O(N__3415),
            .I(un2_r_count_2hz_1_cry_4));
    CascadeMux I__355 (
            .O(N__3412),
            .I(N__3409));
    InMux I__354 (
            .O(N__3409),
            .I(N__3406));
    LocalMux I__353 (
            .O(N__3406),
            .I(o_LED_23_1_and));
    CascadeMux I__352 (
            .O(N__3403),
            .I(N__3400));
    InMux I__351 (
            .O(N__3400),
            .I(N__3397));
    LocalMux I__350 (
            .O(N__3397),
            .I(o_LED_23_0_and));
    CascadeMux I__349 (
            .O(N__3394),
            .I(N__3391));
    InMux I__348 (
            .O(N__3391),
            .I(N__3388));
    LocalMux I__347 (
            .O(N__3388),
            .I(o_LED_23_7_and));
    CascadeMux I__346 (
            .O(N__3385),
            .I(N__3382));
    InMux I__345 (
            .O(N__3382),
            .I(N__3379));
    LocalMux I__344 (
            .O(N__3379),
            .I(o_LED_23_5_and));
    IoInMux I__343 (
            .O(N__3376),
            .I(N__3373));
    LocalMux I__342 (
            .O(N__3373),
            .I(N__3370));
    Span4Mux_s3_h I__341 (
            .O(N__3370),
            .I(N__3366));
    InMux I__340 (
            .O(N__3369),
            .I(N__3363));
    Odrv4 I__339 (
            .O(N__3366),
            .I(o_LED_2_c));
    LocalMux I__338 (
            .O(N__3363),
            .I(o_LED_2_c));
    CascadeMux I__337 (
            .O(N__3358),
            .I(N__3349));
    CascadeMux I__336 (
            .O(N__3357),
            .I(N__3345));
    CascadeMux I__335 (
            .O(N__3356),
            .I(N__3342));
    CascadeMux I__334 (
            .O(N__3355),
            .I(N__3338));
    CascadeMux I__333 (
            .O(N__3354),
            .I(N__3333));
    CascadeMux I__332 (
            .O(N__3353),
            .I(N__3329));
    InMux I__331 (
            .O(N__3352),
            .I(N__3325));
    InMux I__330 (
            .O(N__3349),
            .I(N__3314));
    InMux I__329 (
            .O(N__3348),
            .I(N__3314));
    InMux I__328 (
            .O(N__3345),
            .I(N__3314));
    InMux I__327 (
            .O(N__3342),
            .I(N__3314));
    InMux I__326 (
            .O(N__3341),
            .I(N__3314));
    InMux I__325 (
            .O(N__3338),
            .I(N__3299));
    InMux I__324 (
            .O(N__3337),
            .I(N__3299));
    InMux I__323 (
            .O(N__3336),
            .I(N__3299));
    InMux I__322 (
            .O(N__3333),
            .I(N__3299));
    InMux I__321 (
            .O(N__3332),
            .I(N__3299));
    InMux I__320 (
            .O(N__3329),
            .I(N__3299));
    InMux I__319 (
            .O(N__3328),
            .I(N__3299));
    LocalMux I__318 (
            .O(N__3325),
            .I(o_LED_33_THRU_CO));
    LocalMux I__317 (
            .O(N__3314),
            .I(o_LED_33_THRU_CO));
    LocalMux I__316 (
            .O(N__3299),
            .I(o_LED_33_THRU_CO));
    CascadeMux I__315 (
            .O(N__3292),
            .I(N__3289));
    InMux I__314 (
            .O(N__3289),
            .I(N__3286));
    LocalMux I__313 (
            .O(N__3286),
            .I(N__3283));
    Odrv4 I__312 (
            .O(N__3283),
            .I(o_LED_33_7_and));
    CascadeMux I__311 (
            .O(N__3280),
            .I(N__3277));
    InMux I__310 (
            .O(N__3277),
            .I(N__3274));
    LocalMux I__309 (
            .O(N__3274),
            .I(o_LED_23_2_and));
    CascadeMux I__308 (
            .O(N__3271),
            .I(N__3268));
    InMux I__307 (
            .O(N__3268),
            .I(N__3265));
    LocalMux I__306 (
            .O(N__3265),
            .I(o_LED_23_3_and));
    CascadeMux I__305 (
            .O(N__3262),
            .I(N__3259));
    InMux I__304 (
            .O(N__3259),
            .I(N__3256));
    LocalMux I__303 (
            .O(N__3256),
            .I(o_LED_33_5_and));
    CascadeMux I__302 (
            .O(N__3253),
            .I(N__3250));
    InMux I__301 (
            .O(N__3250),
            .I(N__3247));
    LocalMux I__300 (
            .O(N__3247),
            .I(o_LED_33_0_and));
    CascadeMux I__299 (
            .O(N__3244),
            .I(N__3241));
    InMux I__298 (
            .O(N__3241),
            .I(N__3238));
    LocalMux I__297 (
            .O(N__3238),
            .I(o_LED_33_6_and));
    InMux I__296 (
            .O(N__3235),
            .I(bfn_7_4_0_));
    CascadeMux I__295 (
            .O(N__3232),
            .I(N__3229));
    InMux I__294 (
            .O(N__3229),
            .I(N__3226));
    LocalMux I__293 (
            .O(N__3226),
            .I(o_LED_33_4_and));
    CascadeMux I__292 (
            .O(N__3223),
            .I(N__3220));
    InMux I__291 (
            .O(N__3220),
            .I(N__3217));
    LocalMux I__290 (
            .O(N__3217),
            .I(o_LED_33_3_and));
    InMux I__289 (
            .O(N__3214),
            .I(bfn_6_8_0_));
    CascadeMux I__288 (
            .O(N__3211),
            .I(o_LED_33_THRU_CO_cascade_));
    IoInMux I__287 (
            .O(N__3208),
            .I(N__3205));
    LocalMux I__286 (
            .O(N__3205),
            .I(N__3202));
    Span4Mux_s2_h I__285 (
            .O(N__3202),
            .I(N__3199));
    Span4Mux_h I__284 (
            .O(N__3199),
            .I(N__3195));
    InMux I__283 (
            .O(N__3198),
            .I(N__3192));
    Odrv4 I__282 (
            .O(N__3195),
            .I(o_LED_3_c));
    LocalMux I__281 (
            .O(N__3192),
            .I(o_LED_3_c));
    CascadeMux I__280 (
            .O(N__3187),
            .I(N__3184));
    InMux I__279 (
            .O(N__3184),
            .I(N__3181));
    LocalMux I__278 (
            .O(N__3181),
            .I(o_LED_33_2_and));
    CascadeMux I__277 (
            .O(N__3178),
            .I(N__3175));
    InMux I__276 (
            .O(N__3175),
            .I(N__3172));
    LocalMux I__275 (
            .O(N__3172),
            .I(o_LED_33_1_and));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_9_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_3_0_ (
            .carryinitin(un2_r_count_5hz_1_cry_8),
            .carryinitout(bfn_9_3_0_));
    defparam IN_MUX_bfv_9_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_4_0_ (
            .carryinitin(un2_r_count_5hz_1_cry_16),
            .carryinitout(bfn_9_4_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(un2_r_count_5hz_1_cry_24),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(un2_r_count_2hz_1_cry_8),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(un2_r_count_2hz_1_cry_16),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(un2_r_count_2hz_1_cry_24),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(un2_r_count_1hz_1_cry_8),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(un2_r_count_1hz_1_cry_16),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(un2_r_count_1hz_1_cry_24),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_3_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(un2_r_count_10hz_1_cry_8),
            .carryinitout(bfn_12_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(un2_r_count_10hz_1_cry_16),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(un2_r_count_10hz_1_cry_24),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(o_LED_43),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(o_LED_33),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(o_LED_23),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(o_LED_13),
            .carryinitout(bfn_11_2_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam o_LED_33_0_c_LC_6_7_0.C_ON=1'b1;
    defparam o_LED_33_0_c_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam o_LED_33_0_c_LC_6_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_0_c_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3253),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(o_LED_33_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_1_c_LC_6_7_1.C_ON=1'b1;
    defparam o_LED_33_1_c_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam o_LED_33_1_c_LC_6_7_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_1_c_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3178),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_0),
            .carryout(o_LED_33_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_2_c_LC_6_7_2.C_ON=1'b1;
    defparam o_LED_33_2_c_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam o_LED_33_2_c_LC_6_7_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_2_c_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3187),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_1),
            .carryout(o_LED_33_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_3_c_LC_6_7_3.C_ON=1'b1;
    defparam o_LED_33_3_c_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam o_LED_33_3_c_LC_6_7_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_3_c_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_2),
            .carryout(o_LED_33_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_4_c_LC_6_7_4.C_ON=1'b1;
    defparam o_LED_33_4_c_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam o_LED_33_4_c_LC_6_7_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_4_c_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3232),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_3),
            .carryout(o_LED_33_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_5_c_LC_6_7_5.C_ON=1'b1;
    defparam o_LED_33_5_c_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam o_LED_33_5_c_LC_6_7_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_5_c_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3262),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_4),
            .carryout(o_LED_33_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_6_c_LC_6_7_6.C_ON=1'b1;
    defparam o_LED_33_6_c_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam o_LED_33_6_c_LC_6_7_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_6_c_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3244),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_5),
            .carryout(o_LED_33_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_7_c_LC_6_7_7.C_ON=1'b1;
    defparam o_LED_33_7_c_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam o_LED_33_7_c_LC_6_7_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_33_7_c_LC_6_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3292),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_33_6),
            .carryout(o_LED_33),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_THRU_LUT4_0_LC_6_8_0.C_ON=1'b0;
    defparam o_LED_33_THRU_LUT4_0_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam o_LED_33_THRU_LUT4_0_LC_6_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_LED_33_THRU_LUT4_0_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3214),
            .lcout(o_LED_33_THRU_CO),
            .ltout(o_LED_33_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_17_LC_6_8_1.C_ON=1'b0;
    defparam r_count_2hz_17_LC_6_8_1.SEQ_MODE=4'b1000;
    defparam r_count_2hz_17_LC_6_8_1.LUT_INIT=16'b0000011000000110;
    LogicCell40 r_count_2hz_17_LC_6_8_1 (
            .in0(N__3891),
            .in1(N__3877),
            .in2(N__3211),
            .in3(_gnd_net_),
            .lcout(r_count_2hzZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6484),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LEDZ0Z_3_LC_6_8_4.C_ON=1'b0;
    defparam o_LEDZ0Z_3_LC_6_8_4.SEQ_MODE=4'b1000;
    defparam o_LEDZ0Z_3_LC_6_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 o_LEDZ0Z_3_LC_6_8_4 (
            .in0(_gnd_net_),
            .in1(N__3198),
            .in2(_gnd_net_),
            .in3(N__3352),
            .lcout(o_LED_3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6484),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_2_c_RNO_LC_6_8_5.C_ON=1'b0;
    defparam o_LED_33_2_c_RNO_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam o_LED_33_2_c_RNO_LC_6_8_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_33_2_c_RNO_LC_6_8_5 (
            .in0(N__3863),
            .in1(N__3836),
            .in2(N__4132),
            .in3(N__3806),
            .lcout(o_LED_33_2_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_1_c_RNO_LC_6_8_7.C_ON=1'b0;
    defparam o_LED_33_1_c_RNO_LC_6_8_7.SEQ_MODE=4'b0000;
    defparam o_LED_33_1_c_RNO_LC_6_8_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_33_1_c_RNO_LC_6_8_7 (
            .in0(N__3890),
            .in1(N__3968),
            .in2(N__3634),
            .in3(N__3923),
            .lcout(o_LED_33_1_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_0_c_LC_7_3_0.C_ON=1'b1;
    defparam o_LED_23_0_c_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam o_LED_23_0_c_LC_7_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_0_c_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3403),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(o_LED_23_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_1_c_LC_7_3_1.C_ON=1'b1;
    defparam o_LED_23_1_c_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam o_LED_23_1_c_LC_7_3_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_1_c_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_0),
            .carryout(o_LED_23_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_2_c_LC_7_3_2.C_ON=1'b1;
    defparam o_LED_23_2_c_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam o_LED_23_2_c_LC_7_3_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_2_c_LC_7_3_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3280),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_1),
            .carryout(o_LED_23_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_3_c_LC_7_3_3.C_ON=1'b1;
    defparam o_LED_23_3_c_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam o_LED_23_3_c_LC_7_3_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_3_c_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3271),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_2),
            .carryout(o_LED_23_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_4_c_LC_7_3_4.C_ON=1'b1;
    defparam o_LED_23_4_c_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam o_LED_23_4_c_LC_7_3_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_4_c_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_3),
            .carryout(o_LED_23_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_5_c_LC_7_3_5.C_ON=1'b1;
    defparam o_LED_23_5_c_LC_7_3_5.SEQ_MODE=4'b0000;
    defparam o_LED_23_5_c_LC_7_3_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_5_c_LC_7_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3385),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_4),
            .carryout(o_LED_23_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_6_c_LC_7_3_6.C_ON=1'b1;
    defparam o_LED_23_6_c_LC_7_3_6.SEQ_MODE=4'b0000;
    defparam o_LED_23_6_c_LC_7_3_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_6_c_LC_7_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_5),
            .carryout(o_LED_23_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_7_c_LC_7_3_7.C_ON=1'b1;
    defparam o_LED_23_7_c_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam o_LED_23_7_c_LC_7_3_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_23_7_c_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3394),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_23_6),
            .carryout(o_LED_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_THRU_LUT4_0_LC_7_4_0.C_ON=1'b0;
    defparam o_LED_23_THRU_LUT4_0_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam o_LED_23_THRU_LUT4_0_LC_7_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_LED_23_THRU_LUT4_0_LC_7_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3235),
            .lcout(o_LED_23_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_1_LC_7_6_0.C_ON=1'b0;
    defparam r_count_2hz_1_LC_7_6_0.SEQ_MODE=4'b1000;
    defparam r_count_2hz_1_LC_7_6_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_count_2hz_1_LC_7_6_0 (
            .in0(_gnd_net_),
            .in1(N__3526),
            .in2(_gnd_net_),
            .in3(N__3504),
            .lcout(r_count_2hzZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6488),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_4_c_RNO_LC_7_6_1.C_ON=1'b0;
    defparam o_LED_33_4_c_RNO_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam o_LED_33_4_c_RNO_LC_7_6_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_33_4_c_RNO_LC_7_6_1 (
            .in0(N__3766),
            .in1(N__3427),
            .in2(N__3751),
            .in3(N__3732),
            .lcout(o_LED_33_4_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_10_LC_7_7_0.C_ON=1'b0;
    defparam r_count_2hz_10_LC_7_7_0.SEQ_MODE=4'b1000;
    defparam r_count_2hz_10_LC_7_7_0.LUT_INIT=16'b0000000001011010;
    LogicCell40 r_count_2hz_10_LC_7_7_0 (
            .in0(N__3667),
            .in1(_gnd_net_),
            .in2(N__3691),
            .in3(N__3341),
            .lcout(r_count_2hzZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6487),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_0_LC_7_7_1.C_ON=1'b0;
    defparam r_count_2hz_0_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam r_count_2hz_0_LC_7_7_1.LUT_INIT=16'b0000010100000101;
    LogicCell40 r_count_2hz_0_LC_7_7_1 (
            .in0(N__3525),
            .in1(_gnd_net_),
            .in2(N__3358),
            .in3(_gnd_net_),
            .lcout(r_count_2hzZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6487),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_3_c_RNO_LC_7_7_2.C_ON=1'b0;
    defparam o_LED_33_3_c_RNO_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam o_LED_33_3_c_RNO_LC_7_7_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_33_3_c_RNO_LC_7_7_2 (
            .in0(N__3503),
            .in1(N__3524),
            .in2(N__3484),
            .in3(N__3465),
            .lcout(o_LED_33_3_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_11_LC_7_7_3.C_ON=1'b0;
    defparam r_count_2hz_11_LC_7_7_3.SEQ_MODE=4'b1000;
    defparam r_count_2hz_11_LC_7_7_3.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_2hz_11_LC_7_7_3 (
            .in0(N__3657),
            .in1(_gnd_net_),
            .in2(N__3356),
            .in3(N__3643),
            .lcout(r_count_2hzZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6487),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_9_LC_7_7_4.C_ON=1'b0;
    defparam r_count_2hz_9_LC_7_7_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_9_LC_7_7_4.LUT_INIT=16'b0000000001011010;
    LogicCell40 r_count_2hz_9_LC_7_7_4 (
            .in0(N__3700),
            .in1(_gnd_net_),
            .in2(N__3718),
            .in3(N__3348),
            .lcout(r_count_2hzZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6487),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_5_c_RNO_LC_7_7_5.C_ON=1'b0;
    defparam o_LED_33_5_c_RNO_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam o_LED_33_5_c_RNO_LC_7_7_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_33_5_c_RNO_LC_7_7_5 (
            .in0(N__3604),
            .in1(N__4101),
            .in2(N__3943),
            .in3(N__3780),
            .lcout(o_LED_33_5_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_0_c_RNO_LC_7_7_6.C_ON=1'b0;
    defparam o_LED_33_0_c_RNO_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam o_LED_33_0_c_RNO_LC_7_7_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_33_0_c_RNO_LC_7_7_6 (
            .in0(N__3714),
            .in1(N__3450),
            .in2(N__3690),
            .in3(N__3656),
            .lcout(o_LED_33_0_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_4_LC_7_7_7.C_ON=1'b0;
    defparam r_count_2hz_4_LC_7_7_7.SEQ_MODE=4'b1000;
    defparam r_count_2hz_4_LC_7_7_7.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_2hz_4_LC_7_7_7 (
            .in0(N__3451),
            .in1(_gnd_net_),
            .in2(N__3357),
            .in3(N__3436),
            .lcout(r_count_2hzZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6487),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_16_LC_7_8_0.C_ON=1'b0;
    defparam r_count_2hz_16_LC_7_8_0.SEQ_MODE=4'b1000;
    defparam r_count_2hz_16_LC_7_8_0.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_2hz_16_LC_7_8_0 (
            .in0(N__3907),
            .in1(N__3925),
            .in2(_gnd_net_),
            .in3(N__3332),
            .lcout(r_count_2hzZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_14_LC_7_8_1.C_ON=1'b0;
    defparam r_count_2hz_14_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam r_count_2hz_14_LC_7_8_1.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_2hz_14_LC_7_8_1 (
            .in0(N__3952),
            .in1(_gnd_net_),
            .in2(N__3353),
            .in3(N__3973),
            .lcout(r_count_2hzZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_19_LC_7_8_2.C_ON=1'b0;
    defparam r_count_2hz_19_LC_7_8_2.SEQ_MODE=4'b1000;
    defparam r_count_2hz_19_LC_7_8_2.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_2hz_19_LC_7_8_2 (
            .in0(N__3820),
            .in1(N__3838),
            .in2(_gnd_net_),
            .in3(N__3336),
            .lcout(r_count_2hzZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_6_c_RNO_LC_7_8_3.C_ON=1'b0;
    defparam o_LED_33_6_c_RNO_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam o_LED_33_6_c_RNO_LC_7_8_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_33_6_c_RNO_LC_7_8_3 (
            .in0(N__4054),
            .in1(N__4068),
            .in2(N__4087),
            .in3(N__4035),
            .lcout(o_LED_33_6_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_20_LC_7_8_4.C_ON=1'b0;
    defparam r_count_2hz_20_LC_7_8_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_20_LC_7_8_4.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_2hz_20_LC_7_8_4 (
            .in0(N__3790),
            .in1(N__3808),
            .in2(_gnd_net_),
            .in3(N__3337),
            .lcout(r_count_2hzZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_18_LC_7_8_5.C_ON=1'b0;
    defparam r_count_2hz_18_LC_7_8_5.SEQ_MODE=4'b1000;
    defparam r_count_2hz_18_LC_7_8_5.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_2hz_18_LC_7_8_5 (
            .in0(N__3847),
            .in1(_gnd_net_),
            .in2(N__3354),
            .in3(N__3865),
            .lcout(r_count_2hzZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_12_LC_7_8_6.C_ON=1'b0;
    defparam r_count_2hz_12_LC_7_8_6.SEQ_MODE=4'b1000;
    defparam r_count_2hz_12_LC_7_8_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_2hz_12_LC_7_8_6 (
            .in0(N__3613),
            .in1(N__3633),
            .in2(_gnd_net_),
            .in3(N__3328),
            .lcout(r_count_2hzZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_22_LC_7_8_7.C_ON=1'b0;
    defparam r_count_2hz_22_LC_7_8_7.SEQ_MODE=4'b1000;
    defparam r_count_2hz_22_LC_7_8_7.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_2hz_22_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(N__4111),
            .in2(N__3355),
            .in3(N__4131),
            .lcout(r_count_2hzZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6485),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_33_7_c_RNO_LC_7_9_3.C_ON=1'b0;
    defparam o_LED_33_7_c_RNO_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam o_LED_33_7_c_RNO_LC_7_9_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_33_7_c_RNO_LC_7_9_3 (
            .in0(N__4020),
            .in1(N__4239),
            .in2(N__3991),
            .in3(N__4005),
            .lcout(o_LED_33_7_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_1_LC_8_2_0.C_ON=1'b0;
    defparam r_count_5hz_1_LC_8_2_0.SEQ_MODE=4'b1000;
    defparam r_count_5hz_1_LC_8_2_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_count_5hz_1_LC_8_2_0 (
            .in0(_gnd_net_),
            .in1(N__4185),
            .in2(_gnd_net_),
            .in3(N__4209),
            .lcout(r_count_5hzZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6505),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_2_c_RNO_LC_8_2_4.C_ON=1'b0;
    defparam o_LED_23_2_c_RNO_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam o_LED_23_2_c_RNO_LC_8_2_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_2_c_RNO_LC_8_2_4 (
            .in0(N__4168),
            .in1(N__4184),
            .in2(N__4150),
            .in3(N__4362),
            .lcout(o_LED_23_2_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_3_c_RNO_LC_8_2_5.C_ON=1'b0;
    defparam o_LED_23_3_c_RNO_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam o_LED_23_3_c_RNO_LC_8_2_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_3_c_RNO_LC_8_2_5 (
            .in0(N__4303),
            .in1(N__4288),
            .in2(N__4348),
            .in3(N__4272),
            .lcout(o_LED_23_3_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_0_LC_8_3_0.C_ON=1'b0;
    defparam r_count_5hz_0_LC_8_3_0.SEQ_MODE=4'b1000;
    defparam r_count_5hz_0_LC_8_3_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 r_count_5hz_0_LC_8_3_0 (
            .in0(_gnd_net_),
            .in1(N__4208),
            .in2(_gnd_net_),
            .in3(N__3567),
            .lcout(r_count_5hzZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_7_LC_8_3_1.C_ON=1'b0;
    defparam r_count_5hz_7_LC_8_3_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_7_LC_8_3_1.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_5hz_7_LC_8_3_1 (
            .in0(N__4312),
            .in1(_gnd_net_),
            .in2(N__3571),
            .in3(N__4330),
            .lcout(r_count_5hzZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_12_LC_8_3_2.C_ON=1'b0;
    defparam r_count_5hz_12_LC_8_3_2.SEQ_MODE=4'b1000;
    defparam r_count_5hz_12_LC_8_3_2.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_5hz_12_LC_8_3_2 (
            .in0(N__4572),
            .in1(N__4558),
            .in2(_gnd_net_),
            .in3(N__3558),
            .lcout(r_count_5hzZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_15_LC_8_3_3.C_ON=1'b0;
    defparam r_count_5hz_15_LC_8_3_3.SEQ_MODE=4'b1000;
    defparam r_count_5hz_15_LC_8_3_3.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_5hz_15_LC_8_3_3 (
            .in0(N__4489),
            .in1(_gnd_net_),
            .in2(N__3570),
            .in3(N__4503),
            .lcout(r_count_5hzZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_14_LC_8_3_4.C_ON=1'b0;
    defparam r_count_5hz_14_LC_8_3_4.SEQ_MODE=4'b1000;
    defparam r_count_5hz_14_LC_8_3_4.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_5hz_14_LC_8_3_4 (
            .in0(N__4533),
            .in1(N__4513),
            .in2(_gnd_net_),
            .in3(N__3559),
            .lcout(r_count_5hzZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_1_c_RNO_LC_8_3_5.C_ON=1'b0;
    defparam o_LED_23_1_c_RNO_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam o_LED_23_1_c_RNO_LC_8_3_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 o_LED_23_1_c_RNO_LC_8_3_5 (
            .in0(N__4480),
            .in1(N__4502),
            .in2(N__4210),
            .in3(N__4448),
            .lcout(o_LED_23_1_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_4_LC_8_3_6.C_ON=1'b0;
    defparam r_count_5hz_4_LC_8_3_6.SEQ_MODE=4'b1000;
    defparam r_count_5hz_4_LC_8_3_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_5hz_4_LC_8_3_6 (
            .in0(N__4387),
            .in1(N__4372),
            .in2(_gnd_net_),
            .in3(N__3563),
            .lcout(r_count_5hzZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6501),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_0_c_RNO_LC_8_3_7.C_ON=1'b0;
    defparam o_LED_23_0_c_RNO_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam o_LED_23_0_c_RNO_LC_8_3_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_23_0_c_RNO_LC_8_3_7 (
            .in0(N__4329),
            .in1(N__4386),
            .in2(N__4534),
            .in3(N__4571),
            .lcout(o_LED_23_0_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_7_c_RNO_LC_8_4_0.C_ON=1'b0;
    defparam o_LED_23_7_c_RNO_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam o_LED_23_7_c_RNO_LC_8_4_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_7_c_RNO_LC_8_4_0 (
            .in0(N__4734),
            .in1(N__4752),
            .in2(N__4789),
            .in3(N__4767),
            .lcout(o_LED_23_7_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_16_LC_8_4_1.C_ON=1'b0;
    defparam r_count_5hz_16_LC_8_4_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_16_LC_8_4_1.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_5hz_16_LC_8_4_1 (
            .in0(_gnd_net_),
            .in1(N__4459),
            .in2(N__3568),
            .in3(N__4479),
            .lcout(r_count_5hzZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6497),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_5_c_RNO_LC_8_4_2.C_ON=1'b0;
    defparam o_LED_23_5_c_RNO_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam o_LED_23_5_c_RNO_LC_8_4_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_5_c_RNO_LC_8_4_2 (
            .in0(N__4704),
            .in1(N__4653),
            .in2(N__4672),
            .in3(N__4690),
            .lcout(o_LED_23_5_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LEDZ0Z_2_LC_8_4_3.C_ON=1'b0;
    defparam o_LEDZ0Z_2_LC_8_4_3.SEQ_MODE=4'b1000;
    defparam o_LEDZ0Z_2_LC_8_4_3.LUT_INIT=16'b0000111111110000;
    LogicCell40 o_LEDZ0Z_2_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3569),
            .in3(N__3369),
            .lcout(o_LED_2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6497),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_6_c_RNO_LC_8_4_4.C_ON=1'b0;
    defparam o_LED_23_6_c_RNO_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam o_LED_23_6_c_RNO_LC_8_4_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_6_c_RNO_LC_8_4_4 (
            .in0(N__4635),
            .in1(N__4620),
            .in2(N__4606),
            .in3(N__4587),
            .lcout(o_LED_23_6_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_23_4_c_RNO_LC_8_4_5.C_ON=1'b0;
    defparam o_LED_23_4_c_RNO_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam o_LED_23_4_c_RNO_LC_8_4_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_23_4_c_RNO_LC_8_4_5 (
            .in0(N__4549),
            .in1(N__4258),
            .in2(N__4423),
            .in3(N__4401),
            .lcout(o_LED_23_4_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_17_LC_8_4_6.C_ON=1'b0;
    defparam r_count_5hz_17_LC_8_4_6.SEQ_MODE=4'b1000;
    defparam r_count_5hz_17_LC_8_4_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_5hz_17_LC_8_4_6 (
            .in0(N__4432),
            .in1(N__4450),
            .in2(_gnd_net_),
            .in3(N__3554),
            .lcout(r_count_5hzZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6497),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_1_c_LC_8_6_0.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_1_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_1_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_r_count_2hz_1_cry_1_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__3523),
            .in2(N__3505),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un2_r_count_2hz_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_2_LC_8_6_1.C_ON=1'b1;
    defparam r_count_2hz_2_LC_8_6_1.SEQ_MODE=4'b1000;
    defparam r_count_2hz_2_LC_8_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_2_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__3483),
            .in2(_gnd_net_),
            .in3(N__3469),
            .lcout(r_count_2hzZ0Z_2),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_1),
            .carryout(un2_r_count_2hz_1_cry_2),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_3_LC_8_6_2.C_ON=1'b1;
    defparam r_count_2hz_3_LC_8_6_2.SEQ_MODE=4'b1000;
    defparam r_count_2hz_3_LC_8_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_3_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(N__3466),
            .in2(_gnd_net_),
            .in3(N__3454),
            .lcout(r_count_2hzZ0Z_3),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_2),
            .carryout(un2_r_count_2hz_1_cry_3),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_3_THRU_LUT4_0_LC_8_6_3.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_3_THRU_LUT4_0_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_3_THRU_LUT4_0_LC_8_6_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_3_THRU_LUT4_0_LC_8_6_3 (
            .in0(_gnd_net_),
            .in1(N__3449),
            .in2(_gnd_net_),
            .in3(N__3430),
            .lcout(un2_r_count_2hz_1_cry_3_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_3),
            .carryout(un2_r_count_2hz_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_5_LC_8_6_4.C_ON=1'b1;
    defparam r_count_2hz_5_LC_8_6_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_5_LC_8_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_5_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(N__3426),
            .in2(_gnd_net_),
            .in3(N__3415),
            .lcout(r_count_2hzZ0Z_5),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_4),
            .carryout(un2_r_count_2hz_1_cry_5),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_6_LC_8_6_5.C_ON=1'b1;
    defparam r_count_2hz_6_LC_8_6_5.SEQ_MODE=4'b1000;
    defparam r_count_2hz_6_LC_8_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_6_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(N__3765),
            .in2(_gnd_net_),
            .in3(N__3754),
            .lcout(r_count_2hzZ0Z_6),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_5),
            .carryout(un2_r_count_2hz_1_cry_6),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_7_LC_8_6_6.C_ON=1'b1;
    defparam r_count_2hz_7_LC_8_6_6.SEQ_MODE=4'b1000;
    defparam r_count_2hz_7_LC_8_6_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_7_LC_8_6_6 (
            .in0(_gnd_net_),
            .in1(N__3747),
            .in2(_gnd_net_),
            .in3(N__3736),
            .lcout(r_count_2hzZ0Z_7),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_6),
            .carryout(un2_r_count_2hz_1_cry_7),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_8_LC_8_6_7.C_ON=1'b1;
    defparam r_count_2hz_8_LC_8_6_7.SEQ_MODE=4'b1000;
    defparam r_count_2hz_8_LC_8_6_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_8_LC_8_6_7 (
            .in0(_gnd_net_),
            .in1(N__3733),
            .in2(_gnd_net_),
            .in3(N__3721),
            .lcout(r_count_2hzZ0Z_8),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_7),
            .carryout(un2_r_count_2hz_1_cry_8),
            .clk(N__6492),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_8_THRU_LUT4_0_LC_8_7_0.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_8_THRU_LUT4_0_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_8_THRU_LUT4_0_LC_8_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_8_THRU_LUT4_0_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(N__3713),
            .in2(_gnd_net_),
            .in3(N__3694),
            .lcout(un2_r_count_2hz_1_cry_8_THRU_CO),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(un2_r_count_2hz_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_9_THRU_LUT4_0_LC_8_7_1.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_9_THRU_LUT4_0_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_9_THRU_LUT4_0_LC_8_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_9_THRU_LUT4_0_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(N__3683),
            .in2(_gnd_net_),
            .in3(N__3661),
            .lcout(un2_r_count_2hz_1_cry_9_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_9),
            .carryout(un2_r_count_2hz_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_10_THRU_LUT4_0_LC_8_7_2.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_10_THRU_LUT4_0_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_10_THRU_LUT4_0_LC_8_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_10_THRU_LUT4_0_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__3658),
            .in2(_gnd_net_),
            .in3(N__3637),
            .lcout(un2_r_count_2hz_1_cry_10_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_10),
            .carryout(un2_r_count_2hz_1_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_11_THRU_LUT4_0_LC_8_7_3.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_11_THRU_LUT4_0_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_11_THRU_LUT4_0_LC_8_7_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_11_THRU_LUT4_0_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(N__3632),
            .in2(_gnd_net_),
            .in3(N__3607),
            .lcout(un2_r_count_2hz_1_cry_11_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_11),
            .carryout(un2_r_count_2hz_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_13_LC_8_7_4.C_ON=1'b1;
    defparam r_count_2hz_13_LC_8_7_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_13_LC_8_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_13_LC_8_7_4 (
            .in0(_gnd_net_),
            .in1(N__3603),
            .in2(_gnd_net_),
            .in3(N__3592),
            .lcout(r_count_2hzZ0Z_13),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_12),
            .carryout(un2_r_count_2hz_1_cry_13),
            .clk(N__6489),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_13_THRU_LUT4_0_LC_8_7_5.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_13_THRU_LUT4_0_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_13_THRU_LUT4_0_LC_8_7_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_13_THRU_LUT4_0_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(N__3969),
            .in2(_gnd_net_),
            .in3(N__3946),
            .lcout(un2_r_count_2hz_1_cry_13_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_13),
            .carryout(un2_r_count_2hz_1_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_15_LC_8_7_6.C_ON=1'b1;
    defparam r_count_2hz_15_LC_8_7_6.SEQ_MODE=4'b1000;
    defparam r_count_2hz_15_LC_8_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_15_LC_8_7_6 (
            .in0(_gnd_net_),
            .in1(N__3942),
            .in2(_gnd_net_),
            .in3(N__3928),
            .lcout(r_count_2hzZ0Z_15),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_14),
            .carryout(un2_r_count_2hz_1_cry_15),
            .clk(N__6489),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_15_THRU_LUT4_0_LC_8_7_7.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_15_THRU_LUT4_0_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_15_THRU_LUT4_0_LC_8_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_15_THRU_LUT4_0_LC_8_7_7 (
            .in0(_gnd_net_),
            .in1(N__3924),
            .in2(_gnd_net_),
            .in3(N__3898),
            .lcout(un2_r_count_2hz_1_cry_15_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_15),
            .carryout(un2_r_count_2hz_1_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_16_THRU_LUT4_0_LC_8_8_0.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_16_THRU_LUT4_0_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_16_THRU_LUT4_0_LC_8_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_16_THRU_LUT4_0_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(N__3895),
            .in2(_gnd_net_),
            .in3(N__3868),
            .lcout(un2_r_count_2hz_1_cry_16_THRU_CO),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(un2_r_count_2hz_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_17_THRU_LUT4_0_LC_8_8_1.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_17_THRU_LUT4_0_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_17_THRU_LUT4_0_LC_8_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_17_THRU_LUT4_0_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__3864),
            .in2(_gnd_net_),
            .in3(N__3841),
            .lcout(un2_r_count_2hz_1_cry_17_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_17),
            .carryout(un2_r_count_2hz_1_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_18_THRU_LUT4_0_LC_8_8_2.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_18_THRU_LUT4_0_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_18_THRU_LUT4_0_LC_8_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_18_THRU_LUT4_0_LC_8_8_2 (
            .in0(_gnd_net_),
            .in1(N__3837),
            .in2(_gnd_net_),
            .in3(N__3811),
            .lcout(un2_r_count_2hz_1_cry_18_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_18),
            .carryout(un2_r_count_2hz_1_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_19_THRU_LUT4_0_LC_8_8_3.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_19_THRU_LUT4_0_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_19_THRU_LUT4_0_LC_8_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_19_THRU_LUT4_0_LC_8_8_3 (
            .in0(_gnd_net_),
            .in1(N__3807),
            .in2(_gnd_net_),
            .in3(N__3784),
            .lcout(un2_r_count_2hz_1_cry_19_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_19),
            .carryout(un2_r_count_2hz_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_21_LC_8_8_4.C_ON=1'b1;
    defparam r_count_2hz_21_LC_8_8_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_21_LC_8_8_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_21_LC_8_8_4 (
            .in0(_gnd_net_),
            .in1(N__3781),
            .in2(_gnd_net_),
            .in3(N__3769),
            .lcout(r_count_2hzZ0Z_21),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_20),
            .carryout(un2_r_count_2hz_1_cry_21),
            .clk(N__6486),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_2hz_1_cry_21_THRU_LUT4_0_LC_8_8_5.C_ON=1'b1;
    defparam un2_r_count_2hz_1_cry_21_THRU_LUT4_0_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam un2_r_count_2hz_1_cry_21_THRU_LUT4_0_LC_8_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_2hz_1_cry_21_THRU_LUT4_0_LC_8_8_5 (
            .in0(_gnd_net_),
            .in1(N__4130),
            .in2(_gnd_net_),
            .in3(N__4105),
            .lcout(un2_r_count_2hz_1_cry_21_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_21),
            .carryout(un2_r_count_2hz_1_cry_22),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_23_LC_8_8_6.C_ON=1'b1;
    defparam r_count_2hz_23_LC_8_8_6.SEQ_MODE=4'b1000;
    defparam r_count_2hz_23_LC_8_8_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_23_LC_8_8_6 (
            .in0(_gnd_net_),
            .in1(N__4102),
            .in2(_gnd_net_),
            .in3(N__4090),
            .lcout(r_count_2hzZ0Z_23),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_22),
            .carryout(un2_r_count_2hz_1_cry_23),
            .clk(N__6486),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_24_LC_8_8_7.C_ON=1'b1;
    defparam r_count_2hz_24_LC_8_8_7.SEQ_MODE=4'b1000;
    defparam r_count_2hz_24_LC_8_8_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_24_LC_8_8_7 (
            .in0(_gnd_net_),
            .in1(N__4086),
            .in2(_gnd_net_),
            .in3(N__4072),
            .lcout(r_count_2hzZ0Z_24),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_23),
            .carryout(un2_r_count_2hz_1_cry_24),
            .clk(N__6486),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_25_LC_8_9_0.C_ON=1'b1;
    defparam r_count_2hz_25_LC_8_9_0.SEQ_MODE=4'b1000;
    defparam r_count_2hz_25_LC_8_9_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_25_LC_8_9_0 (
            .in0(_gnd_net_),
            .in1(N__4069),
            .in2(_gnd_net_),
            .in3(N__4057),
            .lcout(r_count_2hzZ0Z_25),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(un2_r_count_2hz_1_cry_25),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_26_LC_8_9_1.C_ON=1'b1;
    defparam r_count_2hz_26_LC_8_9_1.SEQ_MODE=4'b1000;
    defparam r_count_2hz_26_LC_8_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_26_LC_8_9_1 (
            .in0(_gnd_net_),
            .in1(N__4053),
            .in2(_gnd_net_),
            .in3(N__4039),
            .lcout(r_count_2hzZ0Z_26),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_25),
            .carryout(un2_r_count_2hz_1_cry_26),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_27_LC_8_9_2.C_ON=1'b1;
    defparam r_count_2hz_27_LC_8_9_2.SEQ_MODE=4'b1000;
    defparam r_count_2hz_27_LC_8_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_27_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__4036),
            .in2(_gnd_net_),
            .in3(N__4024),
            .lcout(r_count_2hzZ0Z_27),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_26),
            .carryout(un2_r_count_2hz_1_cry_27),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_28_LC_8_9_3.C_ON=1'b1;
    defparam r_count_2hz_28_LC_8_9_3.SEQ_MODE=4'b1000;
    defparam r_count_2hz_28_LC_8_9_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_28_LC_8_9_3 (
            .in0(_gnd_net_),
            .in1(N__4021),
            .in2(_gnd_net_),
            .in3(N__4009),
            .lcout(r_count_2hzZ0Z_28),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_27),
            .carryout(un2_r_count_2hz_1_cry_28),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_29_LC_8_9_4.C_ON=1'b1;
    defparam r_count_2hz_29_LC_8_9_4.SEQ_MODE=4'b1000;
    defparam r_count_2hz_29_LC_8_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_29_LC_8_9_4 (
            .in0(_gnd_net_),
            .in1(N__4006),
            .in2(_gnd_net_),
            .in3(N__3994),
            .lcout(r_count_2hzZ0Z_29),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_28),
            .carryout(un2_r_count_2hz_1_cry_29),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_30_LC_8_9_5.C_ON=1'b1;
    defparam r_count_2hz_30_LC_8_9_5.SEQ_MODE=4'b1000;
    defparam r_count_2hz_30_LC_8_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_2hz_30_LC_8_9_5 (
            .in0(_gnd_net_),
            .in1(N__3990),
            .in2(_gnd_net_),
            .in3(N__3976),
            .lcout(r_count_2hzZ0Z_30),
            .ltout(),
            .carryin(un2_r_count_2hz_1_cry_29),
            .carryout(un2_r_count_2hz_1_cry_30),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_2hz_31_LC_8_9_6.C_ON=1'b0;
    defparam r_count_2hz_31_LC_8_9_6.SEQ_MODE=4'b1000;
    defparam r_count_2hz_31_LC_8_9_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_count_2hz_31_LC_8_9_6 (
            .in0(_gnd_net_),
            .in1(N__4240),
            .in2(_gnd_net_),
            .in3(N__4243),
            .lcout(r_count_2hzZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6490),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_5_LC_8_10_1.C_ON=1'b0;
    defparam r_count_1hz_5_LC_8_10_1.SEQ_MODE=4'b1000;
    defparam r_count_1hz_5_LC_8_10_1.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_5_LC_8_10_1 (
            .in0(N__5001),
            .in1(N__4984),
            .in2(_gnd_net_),
            .in3(N__4868),
            .lcout(r_count_1hzZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6491),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_3_c_RNO_LC_8_10_2.C_ON=1'b0;
    defparam o_LED_43_3_c_RNO_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam o_LED_43_3_c_RNO_LC_8_10_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_43_3_c_RNO_LC_8_10_2 (
            .in0(N__5092),
            .in1(N__5116),
            .in2(N__5065),
            .in3(N__5041),
            .lcout(o_LED_43_3_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LEDZ0Z_4_LC_8_10_4.C_ON=1'b0;
    defparam o_LEDZ0Z_4_LC_8_10_4.SEQ_MODE=4'b1000;
    defparam o_LEDZ0Z_4_LC_8_10_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 o_LEDZ0Z_4_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4876),
            .in3(N__4221),
            .lcout(o_LED_4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6491),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_0_c_RNO_LC_8_10_6.C_ON=1'b0;
    defparam o_LED_43_0_c_RNO_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam o_LED_43_0_c_RNO_LC_8_10_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_43_0_c_RNO_LC_8_10_6 (
            .in0(N__5305),
            .in1(N__5000),
            .in2(N__5269),
            .in3(N__5225),
            .lcout(o_LED_43_0_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_0_LC_8_11_4.C_ON=1'b0;
    defparam r_count_1hz_0_LC_8_11_4.SEQ_MODE=4'b1000;
    defparam r_count_1hz_0_LC_8_11_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 r_count_1hz_0_LC_8_11_4 (
            .in0(_gnd_net_),
            .in1(N__5120),
            .in2(_gnd_net_),
            .in3(N__4872),
            .lcout(r_count_1hzZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6494),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_1_c_LC_9_2_0.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_1_c_LC_9_2_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_1_c_LC_9_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_r_count_5hz_1_cry_1_c_LC_9_2_0 (
            .in0(_gnd_net_),
            .in1(N__4204),
            .in2(N__4186),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(un2_r_count_5hz_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_2_LC_9_2_1.C_ON=1'b1;
    defparam r_count_5hz_2_LC_9_2_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_2_LC_9_2_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_2_LC_9_2_1 (
            .in0(_gnd_net_),
            .in1(N__4164),
            .in2(_gnd_net_),
            .in3(N__4153),
            .lcout(r_count_5hzZ0Z_2),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_1),
            .carryout(un2_r_count_5hz_1_cry_2),
            .clk(N__6509),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_3_LC_9_2_2.C_ON=1'b1;
    defparam r_count_5hz_3_LC_9_2_2.SEQ_MODE=4'b1000;
    defparam r_count_5hz_3_LC_9_2_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_3_LC_9_2_2 (
            .in0(_gnd_net_),
            .in1(N__4146),
            .in2(_gnd_net_),
            .in3(N__4135),
            .lcout(r_count_5hzZ0Z_3),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_2),
            .carryout(un2_r_count_5hz_1_cry_3),
            .clk(N__6509),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_3_THRU_LUT4_0_LC_9_2_3.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_3_THRU_LUT4_0_LC_9_2_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_3_THRU_LUT4_0_LC_9_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_3_THRU_LUT4_0_LC_9_2_3 (
            .in0(_gnd_net_),
            .in1(N__4385),
            .in2(_gnd_net_),
            .in3(N__4366),
            .lcout(un2_r_count_5hz_1_cry_3_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_3),
            .carryout(un2_r_count_5hz_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_5_LC_9_2_4.C_ON=1'b1;
    defparam r_count_5hz_5_LC_9_2_4.SEQ_MODE=4'b1000;
    defparam r_count_5hz_5_LC_9_2_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_5_LC_9_2_4 (
            .in0(_gnd_net_),
            .in1(N__4363),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(r_count_5hzZ0Z_5),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_4),
            .carryout(un2_r_count_5hz_1_cry_5),
            .clk(N__6509),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_6_LC_9_2_5.C_ON=1'b1;
    defparam r_count_5hz_6_LC_9_2_5.SEQ_MODE=4'b1000;
    defparam r_count_5hz_6_LC_9_2_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_6_LC_9_2_5 (
            .in0(_gnd_net_),
            .in1(N__4344),
            .in2(_gnd_net_),
            .in3(N__4333),
            .lcout(r_count_5hzZ0Z_6),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_5),
            .carryout(un2_r_count_5hz_1_cry_6),
            .clk(N__6509),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_6_THRU_LUT4_0_LC_9_2_6.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_6_THRU_LUT4_0_LC_9_2_6.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_6_THRU_LUT4_0_LC_9_2_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_6_THRU_LUT4_0_LC_9_2_6 (
            .in0(_gnd_net_),
            .in1(N__4328),
            .in2(_gnd_net_),
            .in3(N__4306),
            .lcout(un2_r_count_5hz_1_cry_6_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_6),
            .carryout(un2_r_count_5hz_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_8_LC_9_2_7.C_ON=1'b1;
    defparam r_count_5hz_8_LC_9_2_7.SEQ_MODE=4'b1000;
    defparam r_count_5hz_8_LC_9_2_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_8_LC_9_2_7 (
            .in0(_gnd_net_),
            .in1(N__4302),
            .in2(_gnd_net_),
            .in3(N__4291),
            .lcout(r_count_5hzZ0Z_8),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_7),
            .carryout(un2_r_count_5hz_1_cry_8),
            .clk(N__6509),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_9_LC_9_3_0.C_ON=1'b1;
    defparam r_count_5hz_9_LC_9_3_0.SEQ_MODE=4'b1000;
    defparam r_count_5hz_9_LC_9_3_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_9_LC_9_3_0 (
            .in0(_gnd_net_),
            .in1(N__4287),
            .in2(_gnd_net_),
            .in3(N__4276),
            .lcout(r_count_5hzZ0Z_9),
            .ltout(),
            .carryin(bfn_9_3_0_),
            .carryout(un2_r_count_5hz_1_cry_9),
            .clk(N__6506),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_10_LC_9_3_1.C_ON=1'b1;
    defparam r_count_5hz_10_LC_9_3_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_10_LC_9_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_10_LC_9_3_1 (
            .in0(_gnd_net_),
            .in1(N__4273),
            .in2(_gnd_net_),
            .in3(N__4261),
            .lcout(r_count_5hzZ0Z_10),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_9),
            .carryout(un2_r_count_5hz_1_cry_10),
            .clk(N__6506),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_11_LC_9_3_2.C_ON=1'b1;
    defparam r_count_5hz_11_LC_9_3_2.SEQ_MODE=4'b1000;
    defparam r_count_5hz_11_LC_9_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_11_LC_9_3_2 (
            .in0(_gnd_net_),
            .in1(N__4257),
            .in2(_gnd_net_),
            .in3(N__4246),
            .lcout(r_count_5hzZ0Z_11),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_10),
            .carryout(un2_r_count_5hz_1_cry_11),
            .clk(N__6506),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_11_THRU_LUT4_0_LC_9_3_3.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_11_THRU_LUT4_0_LC_9_3_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_11_THRU_LUT4_0_LC_9_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_11_THRU_LUT4_0_LC_9_3_3 (
            .in0(_gnd_net_),
            .in1(N__4573),
            .in2(_gnd_net_),
            .in3(N__4552),
            .lcout(un2_r_count_5hz_1_cry_11_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_11),
            .carryout(un2_r_count_5hz_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_13_LC_9_3_4.C_ON=1'b1;
    defparam r_count_5hz_13_LC_9_3_4.SEQ_MODE=4'b1000;
    defparam r_count_5hz_13_LC_9_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_13_LC_9_3_4 (
            .in0(_gnd_net_),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(N__4537),
            .lcout(r_count_5hzZ0Z_13),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_12),
            .carryout(un2_r_count_5hz_1_cry_13),
            .clk(N__6506),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_13_THRU_LUT4_0_LC_9_3_5.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_13_THRU_LUT4_0_LC_9_3_5.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_13_THRU_LUT4_0_LC_9_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_13_THRU_LUT4_0_LC_9_3_5 (
            .in0(_gnd_net_),
            .in1(N__4532),
            .in2(_gnd_net_),
            .in3(N__4507),
            .lcout(un2_r_count_5hz_1_cry_13_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_13),
            .carryout(un2_r_count_5hz_1_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_14_THRU_LUT4_0_LC_9_3_6.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_14_THRU_LUT4_0_LC_9_3_6.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_14_THRU_LUT4_0_LC_9_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_14_THRU_LUT4_0_LC_9_3_6 (
            .in0(_gnd_net_),
            .in1(N__4504),
            .in2(_gnd_net_),
            .in3(N__4483),
            .lcout(un2_r_count_5hz_1_cry_14_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_14),
            .carryout(un2_r_count_5hz_1_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_15_THRU_LUT4_0_LC_9_3_7.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_15_THRU_LUT4_0_LC_9_3_7.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_15_THRU_LUT4_0_LC_9_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_15_THRU_LUT4_0_LC_9_3_7 (
            .in0(_gnd_net_),
            .in1(N__4478),
            .in2(_gnd_net_),
            .in3(N__4453),
            .lcout(un2_r_count_5hz_1_cry_15_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_15),
            .carryout(un2_r_count_5hz_1_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_5hz_1_cry_16_THRU_LUT4_0_LC_9_4_0.C_ON=1'b1;
    defparam un2_r_count_5hz_1_cry_16_THRU_LUT4_0_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_5hz_1_cry_16_THRU_LUT4_0_LC_9_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_5hz_1_cry_16_THRU_LUT4_0_LC_9_4_0 (
            .in0(_gnd_net_),
            .in1(N__4449),
            .in2(_gnd_net_),
            .in3(N__4426),
            .lcout(un2_r_count_5hz_1_cry_16_THRU_CO),
            .ltout(),
            .carryin(bfn_9_4_0_),
            .carryout(un2_r_count_5hz_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_18_LC_9_4_1.C_ON=1'b1;
    defparam r_count_5hz_18_LC_9_4_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_18_LC_9_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_18_LC_9_4_1 (
            .in0(_gnd_net_),
            .in1(N__4422),
            .in2(_gnd_net_),
            .in3(N__4405),
            .lcout(r_count_5hzZ0Z_18),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_17),
            .carryout(un2_r_count_5hz_1_cry_18),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_19_LC_9_4_2.C_ON=1'b1;
    defparam r_count_5hz_19_LC_9_4_2.SEQ_MODE=4'b1000;
    defparam r_count_5hz_19_LC_9_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_19_LC_9_4_2 (
            .in0(_gnd_net_),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__4390),
            .lcout(r_count_5hzZ0Z_19),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_18),
            .carryout(un2_r_count_5hz_1_cry_19),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_20_LC_9_4_3.C_ON=1'b1;
    defparam r_count_5hz_20_LC_9_4_3.SEQ_MODE=4'b1000;
    defparam r_count_5hz_20_LC_9_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_20_LC_9_4_3 (
            .in0(_gnd_net_),
            .in1(N__4705),
            .in2(_gnd_net_),
            .in3(N__4693),
            .lcout(r_count_5hzZ0Z_20),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_19),
            .carryout(un2_r_count_5hz_1_cry_20),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_21_LC_9_4_4.C_ON=1'b1;
    defparam r_count_5hz_21_LC_9_4_4.SEQ_MODE=4'b1000;
    defparam r_count_5hz_21_LC_9_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_21_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__4675),
            .lcout(r_count_5hzZ0Z_21),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_20),
            .carryout(un2_r_count_5hz_1_cry_21),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_22_LC_9_4_5.C_ON=1'b1;
    defparam r_count_5hz_22_LC_9_4_5.SEQ_MODE=4'b1000;
    defparam r_count_5hz_22_LC_9_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_22_LC_9_4_5 (
            .in0(_gnd_net_),
            .in1(N__4671),
            .in2(_gnd_net_),
            .in3(N__4657),
            .lcout(r_count_5hzZ0Z_22),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_21),
            .carryout(un2_r_count_5hz_1_cry_22),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_23_LC_9_4_6.C_ON=1'b1;
    defparam r_count_5hz_23_LC_9_4_6.SEQ_MODE=4'b1000;
    defparam r_count_5hz_23_LC_9_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_23_LC_9_4_6 (
            .in0(_gnd_net_),
            .in1(N__4654),
            .in2(_gnd_net_),
            .in3(N__4639),
            .lcout(r_count_5hzZ0Z_23),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_22),
            .carryout(un2_r_count_5hz_1_cry_23),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_24_LC_9_4_7.C_ON=1'b1;
    defparam r_count_5hz_24_LC_9_4_7.SEQ_MODE=4'b1000;
    defparam r_count_5hz_24_LC_9_4_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_24_LC_9_4_7 (
            .in0(_gnd_net_),
            .in1(N__4636),
            .in2(_gnd_net_),
            .in3(N__4624),
            .lcout(r_count_5hzZ0Z_24),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_23),
            .carryout(un2_r_count_5hz_1_cry_24),
            .clk(N__6502),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_25_LC_9_5_0.C_ON=1'b1;
    defparam r_count_5hz_25_LC_9_5_0.SEQ_MODE=4'b1000;
    defparam r_count_5hz_25_LC_9_5_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_25_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__4621),
            .in2(_gnd_net_),
            .in3(N__4609),
            .lcout(r_count_5hzZ0Z_25),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(un2_r_count_5hz_1_cry_25),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_26_LC_9_5_1.C_ON=1'b1;
    defparam r_count_5hz_26_LC_9_5_1.SEQ_MODE=4'b1000;
    defparam r_count_5hz_26_LC_9_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_26_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__4605),
            .in2(_gnd_net_),
            .in3(N__4591),
            .lcout(r_count_5hzZ0Z_26),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_25),
            .carryout(un2_r_count_5hz_1_cry_26),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_27_LC_9_5_2.C_ON=1'b1;
    defparam r_count_5hz_27_LC_9_5_2.SEQ_MODE=4'b1000;
    defparam r_count_5hz_27_LC_9_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_27_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(N__4588),
            .in2(_gnd_net_),
            .in3(N__4576),
            .lcout(r_count_5hzZ0Z_27),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_26),
            .carryout(un2_r_count_5hz_1_cry_27),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_28_LC_9_5_3.C_ON=1'b1;
    defparam r_count_5hz_28_LC_9_5_3.SEQ_MODE=4'b1000;
    defparam r_count_5hz_28_LC_9_5_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_28_LC_9_5_3 (
            .in0(_gnd_net_),
            .in1(N__4785),
            .in2(_gnd_net_),
            .in3(N__4771),
            .lcout(r_count_5hzZ0Z_28),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_27),
            .carryout(un2_r_count_5hz_1_cry_28),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_29_LC_9_5_4.C_ON=1'b1;
    defparam r_count_5hz_29_LC_9_5_4.SEQ_MODE=4'b1000;
    defparam r_count_5hz_29_LC_9_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_29_LC_9_5_4 (
            .in0(_gnd_net_),
            .in1(N__4768),
            .in2(_gnd_net_),
            .in3(N__4756),
            .lcout(r_count_5hzZ0Z_29),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_28),
            .carryout(un2_r_count_5hz_1_cry_29),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_30_LC_9_5_5.C_ON=1'b1;
    defparam r_count_5hz_30_LC_9_5_5.SEQ_MODE=4'b1000;
    defparam r_count_5hz_30_LC_9_5_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_5hz_30_LC_9_5_5 (
            .in0(_gnd_net_),
            .in1(N__4753),
            .in2(_gnd_net_),
            .in3(N__4741),
            .lcout(r_count_5hzZ0Z_30),
            .ltout(),
            .carryin(un2_r_count_5hz_1_cry_29),
            .carryout(un2_r_count_5hz_1_cry_30),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_5hz_31_LC_9_5_6.C_ON=1'b0;
    defparam r_count_5hz_31_LC_9_5_6.SEQ_MODE=4'b1000;
    defparam r_count_5hz_31_LC_9_5_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_count_5hz_31_LC_9_5_6 (
            .in0(_gnd_net_),
            .in1(N__4735),
            .in2(_gnd_net_),
            .in3(N__4738),
            .lcout(r_count_5hzZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6499),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_0_c_LC_9_9_0.C_ON=1'b1;
    defparam o_LED_43_0_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam o_LED_43_0_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_0_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4723),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(o_LED_43_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_1_c_LC_9_9_1.C_ON=1'b1;
    defparam o_LED_43_1_c_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam o_LED_43_1_c_LC_9_9_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_1_c_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4807),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_0),
            .carryout(o_LED_43_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_2_c_LC_9_9_2.C_ON=1'b1;
    defparam o_LED_43_2_c_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam o_LED_43_2_c_LC_9_9_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_2_c_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4798),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_1),
            .carryout(o_LED_43_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_3_c_LC_9_9_3.C_ON=1'b1;
    defparam o_LED_43_3_c_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam o_LED_43_3_c_LC_9_9_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_3_c_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4714),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_2),
            .carryout(o_LED_43_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_4_c_LC_9_9_4.C_ON=1'b1;
    defparam o_LED_43_4_c_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam o_LED_43_4_c_LC_9_9_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_4_c_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5143),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_3),
            .carryout(o_LED_43_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_5_c_LC_9_9_5.C_ON=1'b1;
    defparam o_LED_43_5_c_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam o_LED_43_5_c_LC_9_9_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_5_c_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(N__6364),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_4),
            .carryout(o_LED_43_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_6_c_LC_9_9_6.C_ON=1'b1;
    defparam o_LED_43_6_c_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam o_LED_43_6_c_LC_9_9_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_6_c_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_5),
            .carryout(o_LED_43_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_7_c_LC_9_9_7.C_ON=1'b1;
    defparam o_LED_43_7_c_LC_9_9_7.SEQ_MODE=4'b0000;
    defparam o_LED_43_7_c_LC_9_9_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_43_7_c_LC_9_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5740),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_43_6),
            .carryout(o_LED_43),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_THRU_LUT4_0_LC_9_10_0.C_ON=1'b0;
    defparam o_LED_43_THRU_LUT4_0_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam o_LED_43_THRU_LUT4_0_LC_9_10_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_LED_43_THRU_LUT4_0_LC_9_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4813),
            .lcout(o_LED_43_THRU_CO),
            .ltout(o_LED_43_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_15_LC_9_10_1.C_ON=1'b0;
    defparam r_count_1hz_15_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam r_count_1hz_15_LC_9_10_1.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_1hz_15_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(N__5161),
            .in2(N__4810),
            .in3(N__5572),
            .lcout(r_count_1hzZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6495),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_1_c_RNO_LC_9_10_2.C_ON=1'b0;
    defparam o_LED_43_1_c_RNO_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam o_LED_43_1_c_RNO_LC_9_10_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_43_1_c_RNO_LC_9_10_2 (
            .in0(N__5160),
            .in1(N__5192),
            .in2(N__5556),
            .in3(N__5510),
            .lcout(o_LED_43_1_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_10_LC_9_10_3.C_ON=1'b0;
    defparam r_count_1hz_10_LC_9_10_3.SEQ_MODE=4'b1000;
    defparam r_count_1hz_10_LC_9_10_3.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_10_LC_9_10_3 (
            .in0(N__5284),
            .in1(N__5303),
            .in2(_gnd_net_),
            .in3(N__4852),
            .lcout(r_count_1hzZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6495),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_2_c_RNO_LC_9_10_4.C_ON=1'b0;
    defparam o_LED_43_2_c_RNO_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam o_LED_43_2_c_RNO_LC_9_10_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_43_2_c_RNO_LC_9_10_4 (
            .in0(N__5373),
            .in1(N__5441),
            .in2(N__5412),
            .in3(N__5477),
            .lcout(o_LED_43_2_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_12_LC_9_10_5.C_ON=1'b0;
    defparam r_count_1hz_12_LC_9_10_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_12_LC_9_10_5.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_12_LC_9_10_5 (
            .in0(N__5209),
            .in1(N__5229),
            .in2(_gnd_net_),
            .in3(N__4854),
            .lcout(r_count_1hzZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6495),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_13_LC_9_10_6.C_ON=1'b0;
    defparam r_count_1hz_13_LC_9_10_6.SEQ_MODE=4'b1000;
    defparam r_count_1hz_13_LC_9_10_6.LUT_INIT=16'b0000010100001010;
    LogicCell40 r_count_1hz_13_LC_9_10_6 (
            .in0(N__5176),
            .in1(_gnd_net_),
            .in2(N__4873),
            .in3(N__5193),
            .lcout(r_count_1hzZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6495),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_11_LC_9_10_7.C_ON=1'b0;
    defparam r_count_1hz_11_LC_9_10_7.SEQ_MODE=4'b1000;
    defparam r_count_1hz_11_LC_9_10_7.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_11_LC_9_10_7 (
            .in0(N__5245),
            .in1(N__5267),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(r_count_1hzZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6495),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_23_LC_9_11_0.C_ON=1'b0;
    defparam r_count_1hz_23_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam r_count_1hz_23_LC_9_11_0.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_23_LC_9_11_0 (
            .in0(N__5350),
            .in1(N__5372),
            .in2(_gnd_net_),
            .in3(N__4867),
            .lcout(r_count_1hzZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_21_LC_9_11_1.C_ON=1'b0;
    defparam r_count_1hz_21_LC_9_11_1.SEQ_MODE=4'b1000;
    defparam r_count_1hz_21_LC_9_11_1.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_1hz_21_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(N__5389),
            .in2(N__4875),
            .in3(N__5411),
            .lcout(r_count_1hzZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_18_LC_9_11_2.C_ON=1'b0;
    defparam r_count_1hz_18_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam r_count_1hz_18_LC_9_11_2.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_18_LC_9_11_2 (
            .in0(N__5497),
            .in1(N__5518),
            .in2(_gnd_net_),
            .in3(N__4859),
            .lcout(r_count_1hzZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_20_LC_9_11_4.C_ON=1'b0;
    defparam r_count_1hz_20_LC_9_11_4.SEQ_MODE=4'b1000;
    defparam r_count_1hz_20_LC_9_11_4.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_20_LC_9_11_4 (
            .in0(N__5425),
            .in1(N__5445),
            .in2(_gnd_net_),
            .in3(N__4863),
            .lcout(r_count_1hzZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_19_LC_9_11_5.C_ON=1'b0;
    defparam r_count_1hz_19_LC_9_11_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_19_LC_9_11_5.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_1hz_19_LC_9_11_5 (
            .in0(_gnd_net_),
            .in1(N__5461),
            .in2(N__4874),
            .in3(N__5481),
            .lcout(r_count_1hzZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_17_LC_9_11_6.C_ON=1'b0;
    defparam r_count_1hz_17_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam r_count_1hz_17_LC_9_11_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_1hz_17_LC_9_11_6 (
            .in0(N__5533),
            .in1(N__5555),
            .in2(_gnd_net_),
            .in3(N__4858),
            .lcout(r_count_1hzZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6498),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_0_c_LC_11_1_0.C_ON=1'b1;
    defparam o_LED_13_0_c_LC_11_1_0.SEQ_MODE=4'b0000;
    defparam o_LED_13_0_c_LC_11_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_0_c_LC_11_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5677),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(o_LED_13_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_1_c_LC_11_1_1.C_ON=1'b1;
    defparam o_LED_13_1_c_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam o_LED_13_1_c_LC_11_1_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_1_c_LC_11_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4885),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_0),
            .carryout(o_LED_13_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_2_c_LC_11_1_2.C_ON=1'b1;
    defparam o_LED_13_2_c_LC_11_1_2.SEQ_MODE=4'b0000;
    defparam o_LED_13_2_c_LC_11_1_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_2_c_LC_11_1_2 (
            .in0(_gnd_net_),
            .in1(N__5659),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_1),
            .carryout(o_LED_13_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_3_c_LC_11_1_3.C_ON=1'b1;
    defparam o_LED_13_3_c_LC_11_1_3.SEQ_MODE=4'b0000;
    defparam o_LED_13_3_c_LC_11_1_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_3_c_LC_11_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5668),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_2),
            .carryout(o_LED_13_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_4_c_LC_11_1_4.C_ON=1'b1;
    defparam o_LED_13_4_c_LC_11_1_4.SEQ_MODE=4'b0000;
    defparam o_LED_13_4_c_LC_11_1_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_4_c_LC_11_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4936),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_3),
            .carryout(o_LED_13_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_5_c_LC_11_1_5.C_ON=1'b1;
    defparam o_LED_13_5_c_LC_11_1_5.SEQ_MODE=4'b0000;
    defparam o_LED_13_5_c_LC_11_1_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_5_c_LC_11_1_5 (
            .in0(_gnd_net_),
            .in1(N__4924),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_4),
            .carryout(o_LED_13_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_6_c_LC_11_1_6.C_ON=1'b1;
    defparam o_LED_13_6_c_LC_11_1_6.SEQ_MODE=4'b0000;
    defparam o_LED_13_6_c_LC_11_1_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_6_c_LC_11_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_5),
            .carryout(o_LED_13_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_7_c_LC_11_1_7.C_ON=1'b1;
    defparam o_LED_13_7_c_LC_11_1_7.SEQ_MODE=4'b0000;
    defparam o_LED_13_7_c_LC_11_1_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 o_LED_13_7_c_LC_11_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4903),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(o_LED_13_6),
            .carryout(o_LED_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_THRU_LUT4_0_LC_11_2_0.C_ON=1'b0;
    defparam o_LED_13_THRU_LUT4_0_LC_11_2_0.SEQ_MODE=4'b0000;
    defparam o_LED_13_THRU_LUT4_0_LC_11_2_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_LED_13_THRU_LUT4_0_LC_11_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4891),
            .lcout(o_LED_13_THRU_CO),
            .ltout(o_LED_13_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_4_LC_11_2_1.C_ON=1'b0;
    defparam r_count_10hz_4_LC_11_2_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_4_LC_11_2_1.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_10hz_4_LC_11_2_1 (
            .in0(_gnd_net_),
            .in1(N__5911),
            .in2(N__4888),
            .in3(N__5929),
            .lcout(r_count_10hzZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6512),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_1_c_RNO_LC_11_2_7.C_ON=1'b0;
    defparam o_LED_13_1_c_RNO_LC_11_2_7.SEQ_MODE=4'b0000;
    defparam o_LED_13_1_c_RNO_LC_11_2_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_13_1_c_RNO_LC_11_2_7 (
            .in0(N__6035),
            .in1(N__6005),
            .in2(N__6112),
            .in3(N__6263),
            .lcout(o_LED_13_1_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_20_LC_11_3_1.C_ON=1'b0;
    defparam r_count_10hz_20_LC_11_3_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_20_LC_11_3_1.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_10hz_20_LC_11_3_1 (
            .in0(_gnd_net_),
            .in1(N__6247),
            .in2(N__5724),
            .in3(N__6267),
            .lcout(r_count_10hzZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_12_LC_11_3_3.C_ON=1'b0;
    defparam r_count_10hz_12_LC_11_3_3.SEQ_MODE=4'b1000;
    defparam r_count_10hz_12_LC_11_3_3.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_10hz_12_LC_11_3_3 (
            .in0(_gnd_net_),
            .in1(N__6091),
            .in2(N__5721),
            .in3(N__6111),
            .lcout(r_count_10hzZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LEDZ0Z_1_LC_11_3_4.C_ON=1'b0;
    defparam o_LEDZ0Z_1_LC_11_3_4.SEQ_MODE=4'b1000;
    defparam o_LEDZ0Z_1_LC_11_3_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 o_LEDZ0Z_1_LC_11_3_4 (
            .in0(_gnd_net_),
            .in1(N__4947),
            .in2(_gnd_net_),
            .in3(N__5715),
            .lcout(o_LED_1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_17_LC_11_3_5.C_ON=1'b0;
    defparam r_count_10hz_17_LC_11_3_5.SEQ_MODE=4'b1000;
    defparam r_count_10hz_17_LC_11_3_5.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_10hz_17_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(N__5989),
            .in2(N__5723),
            .in3(N__6009),
            .lcout(r_count_10hzZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_9_LC_11_3_6.C_ON=1'b0;
    defparam r_count_10hz_9_LC_11_3_6.SEQ_MODE=4'b1000;
    defparam r_count_10hz_9_LC_11_3_6.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_10hz_9_LC_11_3_6 (
            .in0(N__5800),
            .in1(N__5818),
            .in2(_gnd_net_),
            .in3(N__5714),
            .lcout(r_count_10hzZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_16_LC_11_3_7.C_ON=1'b0;
    defparam r_count_10hz_16_LC_11_3_7.SEQ_MODE=4'b1000;
    defparam r_count_10hz_16_LC_11_3_7.LUT_INIT=16'b0000001100001100;
    LogicCell40 r_count_10hz_16_LC_11_3_7 (
            .in0(_gnd_net_),
            .in1(N__6019),
            .in2(N__5722),
            .in3(N__6037),
            .lcout(r_count_10hzZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6510),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_4_c_RNO_LC_11_4_7.C_ON=1'b0;
    defparam o_LED_13_4_c_RNO_LC_11_4_7.SEQ_MODE=4'b0000;
    defparam o_LED_13_4_c_RNO_LC_11_4_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_4_c_RNO_LC_11_4_7 (
            .in0(N__6051),
            .in1(N__6066),
            .in2(N__5977),
            .in3(N__6081),
            .lcout(o_LED_13_4_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_5_c_RNO_LC_11_5_1.C_ON=1'b0;
    defparam o_LED_13_5_c_RNO_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam o_LED_13_5_c_RNO_LC_11_5_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_5_c_RNO_LC_11_5_1 (
            .in0(N__6195),
            .in1(N__6235),
            .in2(N__6217),
            .in3(N__6285),
            .lcout(o_LED_13_5_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_6_c_RNO_LC_11_5_3.C_ON=1'b0;
    defparam o_LED_13_6_c_RNO_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam o_LED_13_6_c_RNO_LC_11_5_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_6_c_RNO_LC_11_5_3 (
            .in0(N__6180),
            .in1(N__6591),
            .in2(N__6166),
            .in3(N__6147),
            .lcout(o_LED_13_6_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_7_c_RNO_LC_11_5_5.C_ON=1'b0;
    defparam o_LED_13_7_c_RNO_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam o_LED_13_7_c_RNO_LC_11_5_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_7_c_RNO_LC_11_5_5 (
            .in0(N__6543),
            .in1(N__6525),
            .in2(N__6577),
            .in3(N__6558),
            .lcout(o_LED_13_7_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_1_LC_11_8_0.C_ON=1'b0;
    defparam r_count_1hz_1_LC_11_8_0.SEQ_MODE=4'b1000;
    defparam r_count_1hz_1_LC_11_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_count_1hz_1_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(N__5087),
            .in2(_gnd_net_),
            .in3(N__5128),
            .lcout(r_count_1hzZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6493),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_4_c_RNO_LC_11_8_2.C_ON=1'b0;
    defparam o_LED_43_4_c_RNO_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam o_LED_43_4_c_RNO_LC_11_8_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_43_4_c_RNO_LC_11_8_2 (
            .in0(N__4969),
            .in1(N__5020),
            .in2(N__5341),
            .in3(N__5322),
            .lcout(o_LED_43_4_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_1_c_LC_11_9_0.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_1_c_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_1_c_LC_11_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_r_count_1hz_1_cry_1_c_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(N__5127),
            .in2(N__5088),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(un2_r_count_1hz_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_2_LC_11_9_1.C_ON=1'b1;
    defparam r_count_1hz_2_LC_11_9_1.SEQ_MODE=4'b1000;
    defparam r_count_1hz_2_LC_11_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_2_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__5055),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(r_count_1hzZ0Z_2),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_1),
            .carryout(un2_r_count_1hz_1_cry_2),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_3_LC_11_9_2.C_ON=1'b1;
    defparam r_count_1hz_3_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam r_count_1hz_3_LC_11_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_3_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__5037),
            .in2(_gnd_net_),
            .in3(N__5023),
            .lcout(r_count_1hzZ0Z_3),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_2),
            .carryout(un2_r_count_1hz_1_cry_3),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_4_LC_11_9_3.C_ON=1'b1;
    defparam r_count_1hz_4_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam r_count_1hz_4_LC_11_9_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_4_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(N__5019),
            .in2(_gnd_net_),
            .in3(N__5008),
            .lcout(r_count_1hzZ0Z_4),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_3),
            .carryout(un2_r_count_1hz_1_cry_4),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_4_THRU_LUT4_0_LC_11_9_4.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_4_THRU_LUT4_0_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_4_THRU_LUT4_0_LC_11_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_4_THRU_LUT4_0_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__5005),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(un2_r_count_1hz_1_cry_4_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_4),
            .carryout(un2_r_count_1hz_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_6_LC_11_9_5.C_ON=1'b1;
    defparam r_count_1hz_6_LC_11_9_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_6_LC_11_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_6_LC_11_9_5 (
            .in0(_gnd_net_),
            .in1(N__4968),
            .in2(_gnd_net_),
            .in3(N__4957),
            .lcout(r_count_1hzZ0Z_6),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_5),
            .carryout(un2_r_count_1hz_1_cry_6),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_7_LC_11_9_6.C_ON=1'b1;
    defparam r_count_1hz_7_LC_11_9_6.SEQ_MODE=4'b1000;
    defparam r_count_1hz_7_LC_11_9_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_7_LC_11_9_6 (
            .in0(_gnd_net_),
            .in1(N__5337),
            .in2(_gnd_net_),
            .in3(N__5326),
            .lcout(r_count_1hzZ0Z_7),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_6),
            .carryout(un2_r_count_1hz_1_cry_7),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_8_LC_11_9_7.C_ON=1'b1;
    defparam r_count_1hz_8_LC_11_9_7.SEQ_MODE=4'b1000;
    defparam r_count_1hz_8_LC_11_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_8_LC_11_9_7 (
            .in0(_gnd_net_),
            .in1(N__5323),
            .in2(_gnd_net_),
            .in3(N__5311),
            .lcout(r_count_1hzZ0Z_8),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_7),
            .carryout(un2_r_count_1hz_1_cry_8),
            .clk(N__6496),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_9_LC_11_10_0.C_ON=1'b1;
    defparam r_count_1hz_9_LC_11_10_0.SEQ_MODE=4'b1000;
    defparam r_count_1hz_9_LC_11_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_9_LC_11_10_0 (
            .in0(_gnd_net_),
            .in1(N__6390),
            .in2(_gnd_net_),
            .in3(N__5308),
            .lcout(r_count_1hzZ0Z_9),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(un2_r_count_1hz_1_cry_9),
            .clk(N__6500),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_9_THRU_LUT4_0_LC_11_10_1.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_9_THRU_LUT4_0_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_9_THRU_LUT4_0_LC_11_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_9_THRU_LUT4_0_LC_11_10_1 (
            .in0(_gnd_net_),
            .in1(N__5304),
            .in2(_gnd_net_),
            .in3(N__5272),
            .lcout(un2_r_count_1hz_1_cry_9_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_9),
            .carryout(un2_r_count_1hz_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_10_THRU_LUT4_0_LC_11_10_2.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_10_THRU_LUT4_0_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_10_THRU_LUT4_0_LC_11_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_10_THRU_LUT4_0_LC_11_10_2 (
            .in0(_gnd_net_),
            .in1(N__5268),
            .in2(_gnd_net_),
            .in3(N__5233),
            .lcout(un2_r_count_1hz_1_cry_10_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_10),
            .carryout(un2_r_count_1hz_1_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_11_THRU_LUT4_0_LC_11_10_3.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_11_THRU_LUT4_0_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_11_THRU_LUT4_0_LC_11_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_11_THRU_LUT4_0_LC_11_10_3 (
            .in0(_gnd_net_),
            .in1(N__5230),
            .in2(_gnd_net_),
            .in3(N__5197),
            .lcout(un2_r_count_1hz_1_cry_11_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_11),
            .carryout(un2_r_count_1hz_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_12_THRU_LUT4_0_LC_11_10_4.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_12_THRU_LUT4_0_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_12_THRU_LUT4_0_LC_11_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_12_THRU_LUT4_0_LC_11_10_4 (
            .in0(_gnd_net_),
            .in1(N__5194),
            .in2(_gnd_net_),
            .in3(N__5167),
            .lcout(un2_r_count_1hz_1_cry_12_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_12),
            .carryout(un2_r_count_1hz_1_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_14_LC_11_10_5.C_ON=1'b1;
    defparam r_count_1hz_14_LC_11_10_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_14_LC_11_10_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_14_LC_11_10_5 (
            .in0(_gnd_net_),
            .in1(N__6415),
            .in2(_gnd_net_),
            .in3(N__5164),
            .lcout(r_count_1hzZ0Z_14),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_13),
            .carryout(un2_r_count_1hz_1_cry_14),
            .clk(N__6500),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_14_THRU_LUT4_0_LC_11_10_6.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_14_THRU_LUT4_0_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_14_THRU_LUT4_0_LC_11_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_14_THRU_LUT4_0_LC_11_10_6 (
            .in0(_gnd_net_),
            .in1(N__5159),
            .in2(_gnd_net_),
            .in3(N__5563),
            .lcout(un2_r_count_1hz_1_cry_14_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_14),
            .carryout(un2_r_count_1hz_1_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_16_LC_11_10_7.C_ON=1'b1;
    defparam r_count_1hz_16_LC_11_10_7.SEQ_MODE=4'b1000;
    defparam r_count_1hz_16_LC_11_10_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_16_LC_11_10_7 (
            .in0(_gnd_net_),
            .in1(N__6376),
            .in2(_gnd_net_),
            .in3(N__5560),
            .lcout(r_count_1hzZ0Z_16),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_15),
            .carryout(un2_r_count_1hz_1_cry_16),
            .clk(N__6500),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_16_THRU_LUT4_0_LC_11_11_0.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_16_THRU_LUT4_0_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_16_THRU_LUT4_0_LC_11_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_16_THRU_LUT4_0_LC_11_11_0 (
            .in0(_gnd_net_),
            .in1(N__5557),
            .in2(_gnd_net_),
            .in3(N__5521),
            .lcout(un2_r_count_1hz_1_cry_16_THRU_CO),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(un2_r_count_1hz_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_17_THRU_LUT4_0_LC_11_11_1.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_17_THRU_LUT4_0_LC_11_11_1.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_17_THRU_LUT4_0_LC_11_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_17_THRU_LUT4_0_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(N__5517),
            .in2(_gnd_net_),
            .in3(N__5485),
            .lcout(un2_r_count_1hz_1_cry_17_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_17),
            .carryout(un2_r_count_1hz_1_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_18_THRU_LUT4_0_LC_11_11_2.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_18_THRU_LUT4_0_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_18_THRU_LUT4_0_LC_11_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_18_THRU_LUT4_0_LC_11_11_2 (
            .in0(_gnd_net_),
            .in1(N__5482),
            .in2(_gnd_net_),
            .in3(N__5449),
            .lcout(un2_r_count_1hz_1_cry_18_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_18),
            .carryout(un2_r_count_1hz_1_cry_19),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_19_THRU_LUT4_0_LC_11_11_3.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_19_THRU_LUT4_0_LC_11_11_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_19_THRU_LUT4_0_LC_11_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_19_THRU_LUT4_0_LC_11_11_3 (
            .in0(_gnd_net_),
            .in1(N__5446),
            .in2(_gnd_net_),
            .in3(N__5416),
            .lcout(un2_r_count_1hz_1_cry_19_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_19),
            .carryout(un2_r_count_1hz_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_20_THRU_LUT4_0_LC_11_11_4.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_20_THRU_LUT4_0_LC_11_11_4.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_20_THRU_LUT4_0_LC_11_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_20_THRU_LUT4_0_LC_11_11_4 (
            .in0(_gnd_net_),
            .in1(N__5413),
            .in2(_gnd_net_),
            .in3(N__5380),
            .lcout(un2_r_count_1hz_1_cry_20_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_20),
            .carryout(un2_r_count_1hz_1_cry_21),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_22_LC_11_11_5.C_ON=1'b1;
    defparam r_count_1hz_22_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_22_LC_11_11_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_22_LC_11_11_5 (
            .in0(_gnd_net_),
            .in1(N__6403),
            .in2(_gnd_net_),
            .in3(N__5377),
            .lcout(r_count_1hzZ0Z_22),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_21),
            .carryout(un2_r_count_1hz_1_cry_22),
            .clk(N__6503),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_1hz_1_cry_22_THRU_LUT4_0_LC_11_11_6.C_ON=1'b1;
    defparam un2_r_count_1hz_1_cry_22_THRU_LUT4_0_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam un2_r_count_1hz_1_cry_22_THRU_LUT4_0_LC_11_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_1hz_1_cry_22_THRU_LUT4_0_LC_11_11_6 (
            .in0(_gnd_net_),
            .in1(N__5374),
            .in2(_gnd_net_),
            .in3(N__5608),
            .lcout(un2_r_count_1hz_1_cry_22_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_22),
            .carryout(un2_r_count_1hz_1_cry_23),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_24_LC_11_11_7.C_ON=1'b1;
    defparam r_count_1hz_24_LC_11_11_7.SEQ_MODE=4'b1000;
    defparam r_count_1hz_24_LC_11_11_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_24_LC_11_11_7 (
            .in0(_gnd_net_),
            .in1(N__6327),
            .in2(_gnd_net_),
            .in3(N__5605),
            .lcout(r_count_1hzZ0Z_24),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_23),
            .carryout(un2_r_count_1hz_1_cry_24),
            .clk(N__6503),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_25_LC_11_12_0.C_ON=1'b1;
    defparam r_count_1hz_25_LC_11_12_0.SEQ_MODE=4'b1000;
    defparam r_count_1hz_25_LC_11_12_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_25_LC_11_12_0 (
            .in0(_gnd_net_),
            .in1(N__6352),
            .in2(_gnd_net_),
            .in3(N__5602),
            .lcout(r_count_1hzZ0Z_25),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(un2_r_count_1hz_1_cry_25),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_26_LC_11_12_1.C_ON=1'b1;
    defparam r_count_1hz_26_LC_11_12_1.SEQ_MODE=4'b1000;
    defparam r_count_1hz_26_LC_11_12_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_26_LC_11_12_1 (
            .in0(_gnd_net_),
            .in1(N__6340),
            .in2(_gnd_net_),
            .in3(N__5599),
            .lcout(r_count_1hzZ0Z_26),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_25),
            .carryout(un2_r_count_1hz_1_cry_26),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_27_LC_11_12_2.C_ON=1'b1;
    defparam r_count_1hz_27_LC_11_12_2.SEQ_MODE=4'b1000;
    defparam r_count_1hz_27_LC_11_12_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_27_LC_11_12_2 (
            .in0(_gnd_net_),
            .in1(N__6313),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(r_count_1hzZ0Z_27),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_26),
            .carryout(un2_r_count_1hz_1_cry_27),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_28_LC_11_12_3.C_ON=1'b1;
    defparam r_count_1hz_28_LC_11_12_3.SEQ_MODE=4'b1000;
    defparam r_count_1hz_28_LC_11_12_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 r_count_1hz_28_LC_11_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5764),
            .in3(N__5593),
            .lcout(r_count_1hzZ0Z_28),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_27),
            .carryout(un2_r_count_1hz_1_cry_28),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_29_LC_11_12_4.C_ON=1'b1;
    defparam r_count_1hz_29_LC_11_12_4.SEQ_MODE=4'b1000;
    defparam r_count_1hz_29_LC_11_12_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_29_LC_11_12_4 (
            .in0(_gnd_net_),
            .in1(N__5581),
            .in2(_gnd_net_),
            .in3(N__5590),
            .lcout(r_count_1hzZ0Z_29),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_28),
            .carryout(un2_r_count_1hz_1_cry_29),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_30_LC_11_12_5.C_ON=1'b1;
    defparam r_count_1hz_30_LC_11_12_5.SEQ_MODE=4'b1000;
    defparam r_count_1hz_30_LC_11_12_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_1hz_30_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(N__5749),
            .in2(_gnd_net_),
            .in3(N__5587),
            .lcout(r_count_1hzZ0Z_30),
            .ltout(),
            .carryin(un2_r_count_1hz_1_cry_29),
            .carryout(un2_r_count_1hz_1_cry_30),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_1hz_31_LC_11_12_6.C_ON=1'b0;
    defparam r_count_1hz_31_LC_11_12_6.SEQ_MODE=4'b1000;
    defparam r_count_1hz_31_LC_11_12_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 r_count_1hz_31_LC_11_12_6 (
            .in0(N__5773),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5584),
            .lcout(r_count_1hzZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6507),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_7_c_RNO_LC_11_12_7.C_ON=1'b0;
    defparam o_LED_43_7_c_RNO_LC_11_12_7.SEQ_MODE=4'b0000;
    defparam o_LED_43_7_c_RNO_LC_11_12_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_43_7_c_RNO_LC_11_12_7 (
            .in0(N__5580),
            .in1(N__5772),
            .in2(N__5763),
            .in3(N__5748),
            .lcout(o_LED_43_7_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_6_LC_12_2_0.C_ON=1'b0;
    defparam r_count_10hz_6_LC_12_2_0.SEQ_MODE=4'b1000;
    defparam r_count_10hz_6_LC_12_2_0.LUT_INIT=16'b0000000001100110;
    LogicCell40 r_count_10hz_6_LC_12_2_0 (
            .in0(N__5887),
            .in1(N__5869),
            .in2(_gnd_net_),
            .in3(N__5716),
            .lcout(r_count_10hzZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6514),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_7_LC_12_2_1.C_ON=1'b0;
    defparam r_count_10hz_7_LC_12_2_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_7_LC_12_2_1.LUT_INIT=16'b0000011000000110;
    LogicCell40 r_count_10hz_7_LC_12_2_1 (
            .in0(N__5859),
            .in1(N__5842),
            .in2(N__5725),
            .in3(_gnd_net_),
            .lcout(r_count_10hzZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6514),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_0_LC_12_2_2.C_ON=1'b0;
    defparam r_count_10hz_0_LC_12_2_2.SEQ_MODE=4'b1000;
    defparam r_count_10hz_0_LC_12_2_2.LUT_INIT=16'b0000000001010101;
    LogicCell40 r_count_10hz_0_LC_12_2_2 (
            .in0(N__5648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5720),
            .lcout(r_count_10hzZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6514),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_0_c_RNO_LC_12_2_3.C_ON=1'b0;
    defparam o_LED_13_0_c_RNO_LC_12_2_3.SEQ_MODE=4'b0000;
    defparam o_LED_13_0_c_RNO_LC_12_2_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 o_LED_13_0_c_RNO_LC_12_2_3 (
            .in0(N__5886),
            .in1(N__5928),
            .in2(N__5860),
            .in3(N__5816),
            .lcout(o_LED_13_0_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_1_LC_12_2_4.C_ON=1'b0;
    defparam r_count_10hz_1_LC_12_2_4.SEQ_MODE=4'b1000;
    defparam r_count_10hz_1_LC_12_2_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 r_count_10hz_1_LC_12_2_4 (
            .in0(N__5629),
            .in1(_gnd_net_),
            .in2(N__5653),
            .in3(_gnd_net_),
            .lcout(r_count_10hzZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6514),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_3_c_RNO_LC_12_2_5.C_ON=1'b0;
    defparam o_LED_13_3_c_RNO_LC_12_2_5.SEQ_MODE=4'b0000;
    defparam o_LED_13_3_c_RNO_LC_12_2_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_3_c_RNO_LC_12_2_5 (
            .in0(N__5833),
            .in1(N__5902),
            .in2(N__5791),
            .in3(N__6130),
            .lcout(o_LED_13_3_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_13_2_c_RNO_LC_12_2_6.C_ON=1'b0;
    defparam o_LED_13_2_c_RNO_LC_12_2_6.SEQ_MODE=4'b0000;
    defparam o_LED_13_2_c_RNO_LC_12_2_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_13_2_c_RNO_LC_12_2_6 (
            .in0(N__5628),
            .in1(N__5959),
            .in2(N__5652),
            .in3(N__5943),
            .lcout(o_LED_13_2_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_1_c_LC_12_3_0.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_1_c_LC_12_3_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_1_c_LC_12_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un2_r_count_10hz_1_cry_1_c_LC_12_3_0 (
            .in0(_gnd_net_),
            .in1(N__5644),
            .in2(N__5627),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(un2_r_count_10hz_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_2_LC_12_3_1.C_ON=1'b1;
    defparam r_count_10hz_2_LC_12_3_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_2_LC_12_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_2_LC_12_3_1 (
            .in0(_gnd_net_),
            .in1(N__5958),
            .in2(_gnd_net_),
            .in3(N__5947),
            .lcout(r_count_10hzZ0Z_2),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_1),
            .carryout(un2_r_count_10hz_1_cry_2),
            .clk(N__6513),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_3_LC_12_3_2.C_ON=1'b1;
    defparam r_count_10hz_3_LC_12_3_2.SEQ_MODE=4'b1000;
    defparam r_count_10hz_3_LC_12_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_3_LC_12_3_2 (
            .in0(_gnd_net_),
            .in1(N__5944),
            .in2(_gnd_net_),
            .in3(N__5932),
            .lcout(r_count_10hzZ0Z_3),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_2),
            .carryout(un2_r_count_10hz_1_cry_3),
            .clk(N__6513),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_3_THRU_LUT4_0_LC_12_3_3.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_3_THRU_LUT4_0_LC_12_3_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_3_THRU_LUT4_0_LC_12_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_3_THRU_LUT4_0_LC_12_3_3 (
            .in0(_gnd_net_),
            .in1(N__5927),
            .in2(_gnd_net_),
            .in3(N__5905),
            .lcout(un2_r_count_10hz_1_cry_3_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_3),
            .carryout(un2_r_count_10hz_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_5_LC_12_3_4.C_ON=1'b1;
    defparam r_count_10hz_5_LC_12_3_4.SEQ_MODE=4'b1000;
    defparam r_count_10hz_5_LC_12_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_5_LC_12_3_4 (
            .in0(_gnd_net_),
            .in1(N__5901),
            .in2(_gnd_net_),
            .in3(N__5890),
            .lcout(r_count_10hzZ0Z_5),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_4),
            .carryout(un2_r_count_10hz_1_cry_5),
            .clk(N__6513),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_5_THRU_LUT4_0_LC_12_3_5.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_5_THRU_LUT4_0_LC_12_3_5.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_5_THRU_LUT4_0_LC_12_3_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_5_THRU_LUT4_0_LC_12_3_5 (
            .in0(_gnd_net_),
            .in1(N__5885),
            .in2(_gnd_net_),
            .in3(N__5863),
            .lcout(un2_r_count_10hz_1_cry_5_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_5),
            .carryout(un2_r_count_10hz_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_6_THRU_LUT4_0_LC_12_3_6.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_6_THRU_LUT4_0_LC_12_3_6.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_6_THRU_LUT4_0_LC_12_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_6_THRU_LUT4_0_LC_12_3_6 (
            .in0(_gnd_net_),
            .in1(N__5855),
            .in2(_gnd_net_),
            .in3(N__5836),
            .lcout(un2_r_count_10hz_1_cry_6_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_6),
            .carryout(un2_r_count_10hz_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_8_LC_12_3_7.C_ON=1'b1;
    defparam r_count_10hz_8_LC_12_3_7.SEQ_MODE=4'b1000;
    defparam r_count_10hz_8_LC_12_3_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_8_LC_12_3_7 (
            .in0(_gnd_net_),
            .in1(N__5832),
            .in2(_gnd_net_),
            .in3(N__5821),
            .lcout(r_count_10hzZ0Z_8),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_7),
            .carryout(un2_r_count_10hz_1_cry_8),
            .clk(N__6513),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_8_THRU_LUT4_0_LC_12_4_0.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_8_THRU_LUT4_0_LC_12_4_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_8_THRU_LUT4_0_LC_12_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_8_THRU_LUT4_0_LC_12_4_0 (
            .in0(_gnd_net_),
            .in1(N__5817),
            .in2(_gnd_net_),
            .in3(N__5794),
            .lcout(un2_r_count_10hz_1_cry_8_THRU_CO),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(un2_r_count_10hz_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_10_LC_12_4_1.C_ON=1'b1;
    defparam r_count_10hz_10_LC_12_4_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_10_LC_12_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_10_LC_12_4_1 (
            .in0(_gnd_net_),
            .in1(N__5787),
            .in2(_gnd_net_),
            .in3(N__6133),
            .lcout(r_count_10hzZ0Z_10),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_9),
            .carryout(un2_r_count_10hz_1_cry_10),
            .clk(N__6511),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_11_LC_12_4_2.C_ON=1'b1;
    defparam r_count_10hz_11_LC_12_4_2.SEQ_MODE=4'b1000;
    defparam r_count_10hz_11_LC_12_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_11_LC_12_4_2 (
            .in0(_gnd_net_),
            .in1(N__6129),
            .in2(_gnd_net_),
            .in3(N__6115),
            .lcout(r_count_10hzZ0Z_11),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_10),
            .carryout(un2_r_count_10hz_1_cry_11),
            .clk(N__6511),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_11_THRU_LUT4_0_LC_12_4_3.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_11_THRU_LUT4_0_LC_12_4_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_11_THRU_LUT4_0_LC_12_4_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_11_THRU_LUT4_0_LC_12_4_3 (
            .in0(_gnd_net_),
            .in1(N__6110),
            .in2(_gnd_net_),
            .in3(N__6085),
            .lcout(un2_r_count_10hz_1_cry_11_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_11),
            .carryout(un2_r_count_10hz_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_13_LC_12_4_4.C_ON=1'b1;
    defparam r_count_10hz_13_LC_12_4_4.SEQ_MODE=4'b1000;
    defparam r_count_10hz_13_LC_12_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_13_LC_12_4_4 (
            .in0(_gnd_net_),
            .in1(N__6082),
            .in2(_gnd_net_),
            .in3(N__6070),
            .lcout(r_count_10hzZ0Z_13),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_12),
            .carryout(un2_r_count_10hz_1_cry_13),
            .clk(N__6511),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_14_LC_12_4_5.C_ON=1'b1;
    defparam r_count_10hz_14_LC_12_4_5.SEQ_MODE=4'b1000;
    defparam r_count_10hz_14_LC_12_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_14_LC_12_4_5 (
            .in0(_gnd_net_),
            .in1(N__6067),
            .in2(_gnd_net_),
            .in3(N__6055),
            .lcout(r_count_10hzZ0Z_14),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_13),
            .carryout(un2_r_count_10hz_1_cry_14),
            .clk(N__6511),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_15_LC_12_4_6.C_ON=1'b1;
    defparam r_count_10hz_15_LC_12_4_6.SEQ_MODE=4'b1000;
    defparam r_count_10hz_15_LC_12_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_15_LC_12_4_6 (
            .in0(_gnd_net_),
            .in1(N__6052),
            .in2(_gnd_net_),
            .in3(N__6040),
            .lcout(r_count_10hzZ0Z_15),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_14),
            .carryout(un2_r_count_10hz_1_cry_15),
            .clk(N__6511),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_15_THRU_LUT4_0_LC_12_4_7.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_15_THRU_LUT4_0_LC_12_4_7.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_15_THRU_LUT4_0_LC_12_4_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_15_THRU_LUT4_0_LC_12_4_7 (
            .in0(_gnd_net_),
            .in1(N__6036),
            .in2(_gnd_net_),
            .in3(N__6013),
            .lcout(un2_r_count_10hz_1_cry_15_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_15),
            .carryout(un2_r_count_10hz_1_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_16_THRU_LUT4_0_LC_12_5_0.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_16_THRU_LUT4_0_LC_12_5_0.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_16_THRU_LUT4_0_LC_12_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_16_THRU_LUT4_0_LC_12_5_0 (
            .in0(_gnd_net_),
            .in1(N__6010),
            .in2(_gnd_net_),
            .in3(N__5980),
            .lcout(un2_r_count_10hz_1_cry_16_THRU_CO),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(un2_r_count_10hz_1_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_18_LC_12_5_1.C_ON=1'b1;
    defparam r_count_10hz_18_LC_12_5_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_18_LC_12_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_18_LC_12_5_1 (
            .in0(_gnd_net_),
            .in1(N__5976),
            .in2(_gnd_net_),
            .in3(N__5962),
            .lcout(r_count_10hzZ0Z_18),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_17),
            .carryout(un2_r_count_10hz_1_cry_18),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_19_LC_12_5_2.C_ON=1'b1;
    defparam r_count_10hz_19_LC_12_5_2.SEQ_MODE=4'b1000;
    defparam r_count_10hz_19_LC_12_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_19_LC_12_5_2 (
            .in0(_gnd_net_),
            .in1(N__6286),
            .in2(_gnd_net_),
            .in3(N__6271),
            .lcout(r_count_10hzZ0Z_19),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_18),
            .carryout(un2_r_count_10hz_1_cry_19),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam un2_r_count_10hz_1_cry_19_THRU_LUT4_0_LC_12_5_3.C_ON=1'b1;
    defparam un2_r_count_10hz_1_cry_19_THRU_LUT4_0_LC_12_5_3.SEQ_MODE=4'b0000;
    defparam un2_r_count_10hz_1_cry_19_THRU_LUT4_0_LC_12_5_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un2_r_count_10hz_1_cry_19_THRU_LUT4_0_LC_12_5_3 (
            .in0(_gnd_net_),
            .in1(N__6268),
            .in2(_gnd_net_),
            .in3(N__6238),
            .lcout(un2_r_count_10hz_1_cry_19_THRU_CO),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_19),
            .carryout(un2_r_count_10hz_1_cry_20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_21_LC_12_5_4.C_ON=1'b1;
    defparam r_count_10hz_21_LC_12_5_4.SEQ_MODE=4'b1000;
    defparam r_count_10hz_21_LC_12_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_21_LC_12_5_4 (
            .in0(_gnd_net_),
            .in1(N__6234),
            .in2(_gnd_net_),
            .in3(N__6220),
            .lcout(r_count_10hzZ0Z_21),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_20),
            .carryout(un2_r_count_10hz_1_cry_21),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_22_LC_12_5_5.C_ON=1'b1;
    defparam r_count_10hz_22_LC_12_5_5.SEQ_MODE=4'b1000;
    defparam r_count_10hz_22_LC_12_5_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_22_LC_12_5_5 (
            .in0(_gnd_net_),
            .in1(N__6213),
            .in2(_gnd_net_),
            .in3(N__6199),
            .lcout(r_count_10hzZ0Z_22),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_21),
            .carryout(un2_r_count_10hz_1_cry_22),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_23_LC_12_5_6.C_ON=1'b1;
    defparam r_count_10hz_23_LC_12_5_6.SEQ_MODE=4'b1000;
    defparam r_count_10hz_23_LC_12_5_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_23_LC_12_5_6 (
            .in0(_gnd_net_),
            .in1(N__6196),
            .in2(_gnd_net_),
            .in3(N__6184),
            .lcout(r_count_10hzZ0Z_23),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_22),
            .carryout(un2_r_count_10hz_1_cry_23),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_24_LC_12_5_7.C_ON=1'b1;
    defparam r_count_10hz_24_LC_12_5_7.SEQ_MODE=4'b1000;
    defparam r_count_10hz_24_LC_12_5_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_24_LC_12_5_7 (
            .in0(_gnd_net_),
            .in1(N__6181),
            .in2(_gnd_net_),
            .in3(N__6169),
            .lcout(r_count_10hzZ0Z_24),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_23),
            .carryout(un2_r_count_10hz_1_cry_24),
            .clk(N__6508),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_25_LC_12_6_0.C_ON=1'b1;
    defparam r_count_10hz_25_LC_12_6_0.SEQ_MODE=4'b1000;
    defparam r_count_10hz_25_LC_12_6_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_25_LC_12_6_0 (
            .in0(_gnd_net_),
            .in1(N__6165),
            .in2(_gnd_net_),
            .in3(N__6151),
            .lcout(r_count_10hzZ0Z_25),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(un2_r_count_10hz_1_cry_25),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_26_LC_12_6_1.C_ON=1'b1;
    defparam r_count_10hz_26_LC_12_6_1.SEQ_MODE=4'b1000;
    defparam r_count_10hz_26_LC_12_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_26_LC_12_6_1 (
            .in0(_gnd_net_),
            .in1(N__6148),
            .in2(_gnd_net_),
            .in3(N__6136),
            .lcout(r_count_10hzZ0Z_26),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_25),
            .carryout(un2_r_count_10hz_1_cry_26),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_27_LC_12_6_2.C_ON=1'b1;
    defparam r_count_10hz_27_LC_12_6_2.SEQ_MODE=4'b1000;
    defparam r_count_10hz_27_LC_12_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_27_LC_12_6_2 (
            .in0(_gnd_net_),
            .in1(N__6592),
            .in2(_gnd_net_),
            .in3(N__6580),
            .lcout(r_count_10hzZ0Z_27),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_26),
            .carryout(un2_r_count_10hz_1_cry_27),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_28_LC_12_6_3.C_ON=1'b1;
    defparam r_count_10hz_28_LC_12_6_3.SEQ_MODE=4'b1000;
    defparam r_count_10hz_28_LC_12_6_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_28_LC_12_6_3 (
            .in0(_gnd_net_),
            .in1(N__6576),
            .in2(_gnd_net_),
            .in3(N__6562),
            .lcout(r_count_10hzZ0Z_28),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_27),
            .carryout(un2_r_count_10hz_1_cry_28),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_29_LC_12_6_4.C_ON=1'b1;
    defparam r_count_10hz_29_LC_12_6_4.SEQ_MODE=4'b1000;
    defparam r_count_10hz_29_LC_12_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_29_LC_12_6_4 (
            .in0(_gnd_net_),
            .in1(N__6559),
            .in2(_gnd_net_),
            .in3(N__6547),
            .lcout(r_count_10hzZ0Z_29),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_28),
            .carryout(un2_r_count_10hz_1_cry_29),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_30_LC_12_6_5.C_ON=1'b1;
    defparam r_count_10hz_30_LC_12_6_5.SEQ_MODE=4'b1000;
    defparam r_count_10hz_30_LC_12_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 r_count_10hz_30_LC_12_6_5 (
            .in0(_gnd_net_),
            .in1(N__6544),
            .in2(_gnd_net_),
            .in3(N__6532),
            .lcout(r_count_10hzZ0Z_30),
            .ltout(),
            .carryin(un2_r_count_10hz_1_cry_29),
            .carryout(un2_r_count_10hz_1_cry_30),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam r_count_10hz_31_LC_12_6_6.C_ON=1'b0;
    defparam r_count_10hz_31_LC_12_6_6.SEQ_MODE=4'b1000;
    defparam r_count_10hz_31_LC_12_6_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_count_10hz_31_LC_12_6_6 (
            .in0(_gnd_net_),
            .in1(N__6526),
            .in2(_gnd_net_),
            .in3(N__6529),
            .lcout(r_count_10hzZ0Z_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6504),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_5_c_RNO_LC_12_10_1.C_ON=1'b0;
    defparam o_LED_43_5_c_RNO_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam o_LED_43_5_c_RNO_LC_12_10_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_43_5_c_RNO_LC_12_10_1 (
            .in0(N__6414),
            .in1(N__6402),
            .in2(N__6391),
            .in3(N__6375),
            .lcout(o_LED_43_5_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_LED_43_6_c_RNO_LC_12_11_2.C_ON=1'b0;
    defparam o_LED_43_6_c_RNO_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam o_LED_43_6_c_RNO_LC_12_11_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 o_LED_43_6_c_RNO_LC_12_11_2 (
            .in0(N__6351),
            .in1(N__6339),
            .in2(N__6328),
            .in3(N__6312),
            .lcout(o_LED_43_6_and),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // LED_blink
