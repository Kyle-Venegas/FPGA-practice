// make 4 LEDs blink at a rate of 10Hz, 5Hz, 2Hz, 1Hz
module LED_blink
#(
  parameter g_COUNT_10HZ  = 1250000,
  parameter g_COUNT_5HZ   = 250000,
  parameter g_COUNT_2HZ   = 6250000,
  parameter g_COUNT_1HZ   = 

