module VGA_pattern_main (
  input  i_Clk,
  input  i_UART_RX,
  output o_UART_RX,
  )